///////////////////////////////////////////////////////////////////////////////
// vim:set shiftwidth=3 softtabstop=3 expandtab:
// $Id: preprocess 2008-03-13 gac1 $
//
// Module: preprocess.v
// Project: NF2.1
// Description: defines a module for the user data path
//
///////////////////////////////////////////////////////////////////////////////
//Utiliza duas fifos, sendo uma ainterface com módulo anterior e segunda
//empilha cinco primeiras palavras de pacotes TCP
`timescale 1ns/1ps

module simulacao
   #(
      parameter DATA_WIDTH = 64,
      parameter CTRL_WIDTH = DATA_WIDTH/8,
      parameter SRAM_ADDR_WIDTH = 24,
      parameter UDP_REG_SRC_WIDTH = 2
   )
   (
      input  [DATA_WIDTH-1:0]             in_data,
      input  [CTRL_WIDTH-1:0]             in_ctrl,
      input                               in_wr,
      output                              in_rdy,

      output reg [DATA_WIDTH-1:0]         out_data,
      output reg[CTRL_WIDTH-1:0]          out_ctrl,
      output                              out_wr,
      input                               out_rdy,

      // --- Register interface
      input                               reg_req_in,
      input                               reg_ack_in,
      input                               reg_rd_wr_L_in,
      input  [`UDP_REG_ADDR_WIDTH-1:0]    reg_addr_in,
      input  [`CPCI_NF2_DATA_WIDTH-1:0]   reg_data_in,
      input  [UDP_REG_SRC_WIDTH-1:0]      reg_src_in,

      output                              reg_req_out,
      output                              reg_ack_out,
      output                              reg_rd_wr_L_out,
      output  [`UDP_REG_ADDR_WIDTH-1:0]   reg_addr_out,
      output  [`CPCI_NF2_DATA_WIDTH-1:0]  reg_data_out,
      output  [UDP_REG_SRC_WIDTH-1:0]     reg_src_out,

      output reg  [SRAM_ADDR_WIDTH-1:0]   hash_0,
      output reg  [SRAM_ADDR_WIDTH-1:0]   hash_1,
      input                               data_proc,
      input                               ack_proc,
      output reg                          data_pkt,
      output reg                          ack_pkt,

      // misc
      input                                reset,
      input                                clk
   );

   // Define the log2 function
   `LOG2_FUNC

   parameter   CRC_ADDR_WIDTH = 19;
////////////////////////////////////////////////////////////////////////////////
// Copyright (C) 1999-2008 Easics NV.
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//
// Purpose : synthesizable CRC function
//   * polynomial: (0 1 3 4 5 6 7 10 11 14 17 18 23)
//   * data width: 256
//
// Info : tools@easics.be
//        http://www.easics.com
////////////////////////////////////////////////////////////////////////////////

  // polynomial: (0 1 3 4 5 6 7 10 11 14 17 18 23)
  // data width: 256
  // convention: the first serial bit is D[255]
  function [22:0] crcf1;

    input [255:0] Data;
    input [22:0] crc;
    reg [255:0] d;
    reg [22:0] c;
    reg [22:0] newcrc;
  begin
    d = Data;
    c = crc;

    newcrc[0] = d[255] ^ d[254] ^ d[252] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[240] ^ d[239] ^ d[238] ^ d[236] ^ d[235] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[225] ^ d[223] ^ d[222] ^ d[219] ^ d[218] ^ d[217] ^ d[215] ^ d[213] ^ d[211] ^ d[210] ^ d[207] ^ d[206] ^ d[203] ^ d[195] ^ d[194] ^ d[193] ^ d[190] ^ d[189] ^ d[184] ^ d[178] ^ d[176] ^ d[172] ^ d[171] ^ d[168] ^ d[166] ^ d[165] ^ d[162] ^ d[158] ^ d[154] ^ d[152] ^ d[148] ^ d[147] ^ d[144] ^ d[143] ^ d[142] ^ d[140] ^ d[139] ^ d[137] ^ d[136] ^ d[133] ^ d[131] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[119] ^ d[117] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[107] ^ d[104] ^ d[103] ^ d[98] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[81] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[72] ^ d[71] ^ d[68] ^ d[66] ^ d[65] ^ d[62] ^ d[60] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[50] ^ d[49] ^ d[46] ^ d[44] ^ d[43] ^ d[42] ^ d[39] ^ d[38] ^ d[31] ^ d[29] ^ d[26] ^ d[23] ^ d[21] ^ d[18] ^ d[15] ^ d[13] ^ d[10] ^ d[9] ^ d[6] ^ d[5] ^ d[0] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[19] ^ c[21] ^ c[22];
    newcrc[1] = d[254] ^ d[253] ^ d[252] ^ d[250] ^ d[248] ^ d[247] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[238] ^ d[237] ^ d[235] ^ d[233] ^ d[228] ^ d[226] ^ d[225] ^ d[224] ^ d[222] ^ d[220] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[204] ^ d[203] ^ d[196] ^ d[193] ^ d[191] ^ d[189] ^ d[185] ^ d[184] ^ d[179] ^ d[178] ^ d[177] ^ d[176] ^ d[173] ^ d[171] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[163] ^ d[162] ^ d[159] ^ d[158] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[149] ^ d[147] ^ d[145] ^ d[142] ^ d[141] ^ d[139] ^ d[138] ^ d[136] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[130] ^ d[124] ^ d[123] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[116] ^ d[111] ^ d[110] ^ d[107] ^ d[105] ^ d[103] ^ d[99] ^ d[98] ^ d[97] ^ d[92] ^ d[88] ^ d[86] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[80] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[71] ^ d[69] ^ d[68] ^ d[67] ^ d[65] ^ d[63] ^ d[62] ^ d[61] ^ d[55] ^ d[51] ^ d[49] ^ d[47] ^ d[46] ^ d[45] ^ d[42] ^ d[40] ^ d[38] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[27] ^ d[26] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[19] ^ d[18] ^ d[16] ^ d[15] ^ d[14] ^ d[13] ^ d[11] ^ d[9] ^ d[7] ^ d[5] ^ d[1] ^ d[0] ^ c[0] ^ c[2] ^ c[4] ^ c[5] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[14] ^ c[15] ^ c[17] ^ c[19] ^ c[20] ^ c[21];
    newcrc[2] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[239] ^ d[238] ^ d[236] ^ d[234] ^ d[229] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[221] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[205] ^ d[204] ^ d[197] ^ d[194] ^ d[192] ^ d[190] ^ d[186] ^ d[185] ^ d[180] ^ d[179] ^ d[178] ^ d[177] ^ d[174] ^ d[172] ^ d[170] ^ d[169] ^ d[168] ^ d[166] ^ d[164] ^ d[163] ^ d[160] ^ d[159] ^ d[156] ^ d[155] ^ d[154] ^ d[153] ^ d[150] ^ d[148] ^ d[146] ^ d[143] ^ d[142] ^ d[140] ^ d[139] ^ d[137] ^ d[135] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[112] ^ d[111] ^ d[108] ^ d[106] ^ d[104] ^ d[100] ^ d[99] ^ d[98] ^ d[93] ^ d[89] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[72] ^ d[70] ^ d[69] ^ d[68] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[56] ^ d[52] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[43] ^ d[41] ^ d[39] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[28] ^ d[27] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[20] ^ d[19] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[12] ^ d[10] ^ d[8] ^ d[6] ^ d[2] ^ d[1] ^ c[1] ^ c[3] ^ c[5] ^ c[6] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[18] ^ c[20] ^ c[21] ^ c[22];
    newcrc[3] = d[250] ^ d[248] ^ d[247] ^ d[245] ^ d[244] ^ d[242] ^ d[238] ^ d[237] ^ d[236] ^ d[232] ^ d[231] ^ d[229] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[216] ^ d[214] ^ d[213] ^ d[212] ^ d[211] ^ d[208] ^ d[207] ^ d[205] ^ d[203] ^ d[198] ^ d[194] ^ d[191] ^ d[190] ^ d[189] ^ d[187] ^ d[186] ^ d[184] ^ d[181] ^ d[180] ^ d[179] ^ d[176] ^ d[175] ^ d[173] ^ d[172] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[166] ^ d[164] ^ d[162] ^ d[161] ^ d[160] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[152] ^ d[151] ^ d[149] ^ d[148] ^ d[142] ^ d[141] ^ d[139] ^ d[138] ^ d[137] ^ d[135] ^ d[134] ^ d[132] ^ d[131] ^ d[129] ^ d[128] ^ d[127] ^ d[124] ^ d[123] ^ d[120] ^ d[118] ^ d[117] ^ d[115] ^ d[114] ^ d[111] ^ d[108] ^ d[105] ^ d[104] ^ d[103] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[96] ^ d[95] ^ d[93] ^ d[92] ^ d[90] ^ d[88] ^ d[86] ^ d[85] ^ d[82] ^ d[81] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[53] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[43] ^ d[40] ^ d[39] ^ d[38] ^ d[34] ^ d[33] ^ d[32] ^ d[28] ^ d[25] ^ d[24] ^ d[20] ^ d[17] ^ d[16] ^ d[11] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[3] ^ d[2] ^ d[0] ^ c[3] ^ c[4] ^ c[5] ^ c[9] ^ c[11] ^ c[12] ^ c[14] ^ c[15] ^ c[17];
    newcrc[4] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[242] ^ d[240] ^ d[237] ^ d[236] ^ d[235] ^ d[233] ^ d[231] ^ d[229] ^ d[227] ^ d[226] ^ d[224] ^ d[223] ^ d[222] ^ d[219] ^ d[218] ^ d[214] ^ d[212] ^ d[211] ^ d[210] ^ d[209] ^ d[208] ^ d[207] ^ d[204] ^ d[203] ^ d[199] ^ d[194] ^ d[193] ^ d[192] ^ d[191] ^ d[189] ^ d[188] ^ d[187] ^ d[185] ^ d[184] ^ d[182] ^ d[181] ^ d[180] ^ d[178] ^ d[177] ^ d[174] ^ d[173] ^ d[172] ^ d[170] ^ d[169] ^ d[167] ^ d[166] ^ d[163] ^ d[161] ^ d[159] ^ d[157] ^ d[156] ^ d[154] ^ d[153] ^ d[150] ^ d[149] ^ d[148] ^ d[147] ^ d[144] ^ d[138] ^ d[137] ^ d[135] ^ d[132] ^ d[131] ^ d[130] ^ d[127] ^ d[126] ^ d[122] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[113] ^ d[111] ^ d[108] ^ d[107] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[95] ^ d[92] ^ d[91] ^ d[89] ^ d[84] ^ d[82] ^ d[81] ^ d[79] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[58] ^ d[55] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[43] ^ d[42] ^ d[41] ^ d[40] ^ d[38] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[25] ^ d[23] ^ d[17] ^ d[15] ^ d[13] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[7] ^ d[5] ^ d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[0] ^ c[2] ^ c[3] ^ c[4] ^ c[7] ^ c[9] ^ c[18] ^ c[19] ^ c[21] ^ c[22];
    newcrc[5] = d[254] ^ d[253] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[237] ^ d[235] ^ d[234] ^ d[231] ^ d[229] ^ d[227] ^ d[224] ^ d[222] ^ d[220] ^ d[218] ^ d[217] ^ d[212] ^ d[209] ^ d[208] ^ d[207] ^ d[206] ^ d[205] ^ d[204] ^ d[203] ^ d[200] ^ d[192] ^ d[188] ^ d[186] ^ d[185] ^ d[184] ^ d[183] ^ d[182] ^ d[181] ^ d[179] ^ d[176] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[170] ^ d[167] ^ d[166] ^ d[165] ^ d[164] ^ d[160] ^ d[157] ^ d[155] ^ d[152] ^ d[151] ^ d[150] ^ d[149] ^ d[147] ^ d[145] ^ d[144] ^ d[143] ^ d[142] ^ d[140] ^ d[138] ^ d[137] ^ d[132] ^ d[129] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[118] ^ d[113] ^ d[111] ^ d[106] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[95] ^ d[94] ^ d[90] ^ d[87] ^ d[86] ^ d[85] ^ d[84] ^ d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[73] ^ d[72] ^ d[70] ^ d[67] ^ d[66] ^ d[64] ^ d[63] ^ d[60] ^ d[58] ^ d[57] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[41] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[32] ^ d[31] ^ d[29] ^ d[24] ^ d[23] ^ d[21] ^ d[16] ^ d[15] ^ d[14] ^ d[12] ^ d[11] ^ d[8] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[1] ^ c[2] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[20] ^ c[21];
    newcrc[6] = d[252] ^ d[250] ^ d[248] ^ d[247] ^ d[245] ^ d[241] ^ d[239] ^ d[231] ^ d[229] ^ d[222] ^ d[221] ^ d[217] ^ d[215] ^ d[211] ^ d[209] ^ d[208] ^ d[205] ^ d[204] ^ d[203] ^ d[201] ^ d[195] ^ d[194] ^ d[190] ^ d[187] ^ d[186] ^ d[185] ^ d[183] ^ d[182] ^ d[180] ^ d[178] ^ d[177] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[167] ^ d[162] ^ d[161] ^ d[156] ^ d[154] ^ d[153] ^ d[151] ^ d[150] ^ d[147] ^ d[146] ^ d[145] ^ d[142] ^ d[141] ^ d[140] ^ d[138] ^ d[137] ^ d[136] ^ d[131] ^ d[130] ^ d[129] ^ d[128] ^ d[123] ^ d[121] ^ d[117] ^ d[115] ^ d[113] ^ d[111] ^ d[109] ^ d[108] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[98] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[88] ^ d[85] ^ d[84] ^ d[82] ^ d[80] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[72] ^ d[67] ^ d[66] ^ d[64] ^ d[62] ^ d[61] ^ d[60] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[18] ^ d[17] ^ d[16] ^ d[12] ^ d[10] ^ d[6] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[6] ^ c[8] ^ c[12] ^ c[14] ^ c[15] ^ c[17] ^ c[19];
    newcrc[7] = d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[251] ^ d[245] ^ d[243] ^ d[239] ^ d[238] ^ d[236] ^ d[235] ^ d[231] ^ d[229] ^ d[228] ^ d[225] ^ d[219] ^ d[217] ^ d[216] ^ d[215] ^ d[213] ^ d[212] ^ d[211] ^ d[209] ^ d[207] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[196] ^ d[194] ^ d[193] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[186] ^ d[183] ^ d[181] ^ d[179] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[166] ^ d[165] ^ d[163] ^ d[158] ^ d[157] ^ d[155] ^ d[151] ^ d[146] ^ d[144] ^ d[141] ^ d[140] ^ d[138] ^ d[136] ^ d[133] ^ d[132] ^ d[130] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[121] ^ d[119] ^ d[118] ^ d[117] ^ d[116] ^ d[115] ^ d[113] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[89] ^ d[87] ^ d[85] ^ d[84] ^ d[79] ^ d[76] ^ d[75] ^ d[73] ^ d[72] ^ d[71] ^ d[67] ^ d[66] ^ d[63] ^ d[61] ^ d[60] ^ d[59] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[37] ^ d[36] ^ d[34] ^ d[33] ^ d[32] ^ d[30] ^ d[29] ^ d[27] ^ d[25] ^ d[24] ^ d[22] ^ d[21] ^ d[19] ^ d[17] ^ d[15] ^ d[11] ^ d[10] ^ d[9] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[10] ^ c[12] ^ c[18] ^ c[19] ^ c[20] ^ c[21] ^ c[22];
    newcrc[8] = d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[246] ^ d[244] ^ d[240] ^ d[239] ^ d[237] ^ d[236] ^ d[232] ^ d[230] ^ d[229] ^ d[226] ^ d[220] ^ d[218] ^ d[217] ^ d[216] ^ d[214] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[205] ^ d[204] ^ d[203] ^ d[197] ^ d[195] ^ d[194] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[184] ^ d[182] ^ d[180] ^ d[176] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[167] ^ d[166] ^ d[164] ^ d[159] ^ d[158] ^ d[156] ^ d[152] ^ d[147] ^ d[145] ^ d[142] ^ d[141] ^ d[139] ^ d[137] ^ d[134] ^ d[133] ^ d[131] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[122] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[112] ^ d[111] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[100] ^ d[99] ^ d[97] ^ d[90] ^ d[88] ^ d[86] ^ d[85] ^ d[80] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[68] ^ d[67] ^ d[64] ^ d[62] ^ d[61] ^ d[60] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[38] ^ d[37] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[30] ^ d[28] ^ d[26] ^ d[25] ^ d[23] ^ d[22] ^ d[20] ^ d[18] ^ d[16] ^ d[12] ^ d[11] ^ d[10] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[11] ^ c[13] ^ c[19] ^ c[20] ^ c[21] ^ c[22];
    newcrc[9] = d[255] ^ d[254] ^ d[253] ^ d[247] ^ d[245] ^ d[241] ^ d[240] ^ d[238] ^ d[237] ^ d[233] ^ d[231] ^ d[230] ^ d[227] ^ d[221] ^ d[219] ^ d[218] ^ d[217] ^ d[215] ^ d[214] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[206] ^ d[205] ^ d[204] ^ d[198] ^ d[196] ^ d[195] ^ d[193] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[185] ^ d[183] ^ d[181] ^ d[177] ^ d[176] ^ d[175] ^ d[174] ^ d[173] ^ d[168] ^ d[167] ^ d[165] ^ d[160] ^ d[159] ^ d[157] ^ d[153] ^ d[148] ^ d[146] ^ d[143] ^ d[142] ^ d[140] ^ d[138] ^ d[135] ^ d[134] ^ d[132] ^ d[130] ^ d[129] ^ d[128] ^ d[127] ^ d[123] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[117] ^ d[115] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[101] ^ d[100] ^ d[98] ^ d[91] ^ d[89] ^ d[87] ^ d[86] ^ d[81] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[69] ^ d[68] ^ d[65] ^ d[63] ^ d[62] ^ d[61] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[50] ^ d[49] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[39] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[32] ^ d[31] ^ d[29] ^ d[27] ^ d[26] ^ d[24] ^ d[23] ^ d[21] ^ d[19] ^ d[17] ^ d[13] ^ d[12] ^ d[11] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[2] ^ c[0] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[12] ^ c[14] ^ c[20] ^ c[21] ^ c[22];
    newcrc[10] = d[252] ^ d[249] ^ d[245] ^ d[243] ^ d[241] ^ d[240] ^ d[236] ^ d[235] ^ d[234] ^ d[230] ^ d[229] ^ d[225] ^ d[223] ^ d[220] ^ d[217] ^ d[216] ^ d[214] ^ d[213] ^ d[212] ^ d[211] ^ d[208] ^ d[205] ^ d[203] ^ d[199] ^ d[197] ^ d[196] ^ d[195] ^ d[192] ^ d[191] ^ d[186] ^ d[182] ^ d[177] ^ d[175] ^ d[174] ^ d[172] ^ d[171] ^ d[169] ^ d[165] ^ d[162] ^ d[161] ^ d[160] ^ d[152] ^ d[149] ^ d[148] ^ d[142] ^ d[141] ^ d[140] ^ d[137] ^ d[135] ^ d[130] ^ d[127] ^ d[126] ^ d[125] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[115] ^ d[112] ^ d[110] ^ d[109] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[95] ^ d[94] ^ d[93] ^ d[90] ^ d[88] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[81] ^ d[77] ^ d[76] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[65] ^ d[64] ^ d[63] ^ d[60] ^ d[59] ^ d[58] ^ d[54] ^ d[53] ^ d[51] ^ d[48] ^ d[45] ^ d[44] ^ d[43] ^ d[42] ^ d[40] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[33] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[15] ^ d[14] ^ d[12] ^ d[8] ^ d[7] ^ d[4] ^ d[3] ^ d[0] ^ c[1] ^ c[2] ^ c[3] ^ c[7] ^ c[8] ^ c[10] ^ c[12] ^ c[16] ^ c[19];
    newcrc[11] = d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[250] ^ d[249] ^ d[248] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[237] ^ d[232] ^ d[229] ^ d[228] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[221] ^ d[219] ^ d[214] ^ d[212] ^ d[211] ^ d[210] ^ d[209] ^ d[207] ^ d[204] ^ d[203] ^ d[200] ^ d[198] ^ d[197] ^ d[196] ^ d[195] ^ d[194] ^ d[192] ^ d[190] ^ d[189] ^ d[187] ^ d[184] ^ d[183] ^ d[175] ^ d[173] ^ d[171] ^ d[170] ^ d[168] ^ d[165] ^ d[163] ^ d[161] ^ d[158] ^ d[154] ^ d[153] ^ d[152] ^ d[150] ^ d[149] ^ d[148] ^ d[147] ^ d[144] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[133] ^ d[129] ^ d[125] ^ d[124] ^ d[122] ^ d[118] ^ d[116] ^ d[115] ^ d[114] ^ d[112] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[102] ^ d[100] ^ d[99] ^ d[98] ^ d[97] ^ d[93] ^ d[92] ^ d[91] ^ d[89] ^ d[86] ^ d[85] ^ d[82] ^ d[81] ^ d[79] ^ d[75] ^ d[74] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[64] ^ d[62] ^ d[61] ^ d[58] ^ d[57] ^ d[56] ^ d[54] ^ d[52] ^ d[50] ^ d[45] ^ d[42] ^ d[41] ^ d[37] ^ d[36] ^ d[34] ^ d[33] ^ d[32] ^ d[30] ^ d[28] ^ d[27] ^ d[25] ^ d[24] ^ d[22] ^ d[18] ^ d[16] ^ d[10] ^ d[8] ^ d[6] ^ d[4] ^ d[1] ^ d[0] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[12] ^ c[15] ^ c[16] ^ c[17] ^ c[19] ^ c[20] ^ c[21] ^ c[22];
    newcrc[12] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[249] ^ d[246] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[233] ^ d[230] ^ d[229] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[215] ^ d[213] ^ d[212] ^ d[211] ^ d[210] ^ d[208] ^ d[205] ^ d[204] ^ d[201] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[195] ^ d[193] ^ d[191] ^ d[190] ^ d[188] ^ d[185] ^ d[184] ^ d[176] ^ d[174] ^ d[172] ^ d[171] ^ d[169] ^ d[166] ^ d[164] ^ d[162] ^ d[159] ^ d[155] ^ d[154] ^ d[153] ^ d[151] ^ d[150] ^ d[149] ^ d[148] ^ d[145] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[134] ^ d[130] ^ d[126] ^ d[125] ^ d[123] ^ d[119] ^ d[117] ^ d[116] ^ d[115] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[103] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[94] ^ d[93] ^ d[92] ^ d[90] ^ d[87] ^ d[86] ^ d[83] ^ d[82] ^ d[80] ^ d[76] ^ d[75] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[65] ^ d[63] ^ d[62] ^ d[59] ^ d[58] ^ d[57] ^ d[55] ^ d[53] ^ d[51] ^ d[46] ^ d[43] ^ d[42] ^ d[38] ^ d[37] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[29] ^ d[28] ^ d[26] ^ d[25] ^ d[23] ^ d[19] ^ d[17] ^ d[11] ^ d[9] ^ d[7] ^ d[5] ^ d[2] ^ d[1] ^ c[0] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[13] ^ c[16] ^ c[17] ^ c[18] ^ c[20] ^ c[21] ^ c[22];
    newcrc[13] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[250] ^ d[247] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[234] ^ d[231] ^ d[230] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[221] ^ d[216] ^ d[214] ^ d[213] ^ d[212] ^ d[211] ^ d[209] ^ d[206] ^ d[205] ^ d[202] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[194] ^ d[192] ^ d[191] ^ d[189] ^ d[186] ^ d[185] ^ d[177] ^ d[175] ^ d[173] ^ d[172] ^ d[170] ^ d[167] ^ d[165] ^ d[163] ^ d[160] ^ d[156] ^ d[155] ^ d[154] ^ d[152] ^ d[151] ^ d[150] ^ d[149] ^ d[146] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[135] ^ d[131] ^ d[127] ^ d[126] ^ d[124] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[114] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[95] ^ d[94] ^ d[93] ^ d[91] ^ d[88] ^ d[87] ^ d[84] ^ d[83] ^ d[81] ^ d[77] ^ d[76] ^ d[75] ^ d[72] ^ d[71] ^ d[70] ^ d[66] ^ d[64] ^ d[63] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[54] ^ d[52] ^ d[47] ^ d[44] ^ d[43] ^ d[39] ^ d[38] ^ d[36] ^ d[35] ^ d[34] ^ d[32] ^ d[30] ^ d[29] ^ d[27] ^ d[26] ^ d[24] ^ d[20] ^ d[18] ^ d[12] ^ d[10] ^ d[8] ^ d[6] ^ d[3] ^ d[2] ^ c[1] ^ c[6] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[14] ^ c[17] ^ c[18] ^ c[19] ^ c[21] ^ c[22];
    newcrc[14] = d[254] ^ d[253] ^ d[251] ^ d[249] ^ d[247] ^ d[245] ^ d[244] ^ d[241] ^ d[239] ^ d[238] ^ d[236] ^ d[230] ^ d[227] ^ d[226] ^ d[224] ^ d[223] ^ d[219] ^ d[218] ^ d[214] ^ d[212] ^ d[211] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[194] ^ d[192] ^ d[189] ^ d[187] ^ d[186] ^ d[184] ^ d[174] ^ d[173] ^ d[172] ^ d[165] ^ d[164] ^ d[162] ^ d[161] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[154] ^ d[153] ^ d[151] ^ d[150] ^ d[148] ^ d[141] ^ d[139] ^ d[137] ^ d[133] ^ d[132] ^ d[131] ^ d[129] ^ d[126] ^ d[124] ^ d[122] ^ d[118] ^ d[114] ^ d[110] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[98] ^ d[93] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[79] ^ d[76] ^ d[75] ^ d[74] ^ d[73] ^ d[68] ^ d[67] ^ d[66] ^ d[64] ^ d[62] ^ d[61] ^ d[58] ^ d[56] ^ d[53] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[40] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[33] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[23] ^ d[19] ^ d[18] ^ d[15] ^ d[11] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[3] ^ d[0] ^ c[3] ^ c[5] ^ c[6] ^ c[8] ^ c[11] ^ c[12] ^ c[14] ^ c[16] ^ c[18] ^ c[20] ^ c[21];
    newcrc[15] = d[255] ^ d[254] ^ d[252] ^ d[250] ^ d[248] ^ d[246] ^ d[245] ^ d[242] ^ d[240] ^ d[239] ^ d[237] ^ d[231] ^ d[228] ^ d[227] ^ d[225] ^ d[224] ^ d[220] ^ d[219] ^ d[215] ^ d[213] ^ d[212] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[195] ^ d[193] ^ d[190] ^ d[188] ^ d[187] ^ d[185] ^ d[175] ^ d[174] ^ d[173] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[159] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[154] ^ d[152] ^ d[151] ^ d[149] ^ d[142] ^ d[140] ^ d[138] ^ d[134] ^ d[133] ^ d[132] ^ d[130] ^ d[127] ^ d[125] ^ d[123] ^ d[119] ^ d[115] ^ d[111] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[103] ^ d[102] ^ d[101] ^ d[99] ^ d[94] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[84] ^ d[83] ^ d[82] ^ d[80] ^ d[77] ^ d[76] ^ d[75] ^ d[74] ^ d[69] ^ d[68] ^ d[67] ^ d[65] ^ d[63] ^ d[62] ^ d[59] ^ d[57] ^ d[54] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[46] ^ d[44] ^ d[43] ^ d[41] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[34] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[24] ^ d[20] ^ d[19] ^ d[16] ^ d[12] ^ d[11] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[1] ^ c[4] ^ c[6] ^ c[7] ^ c[9] ^ c[12] ^ c[13] ^ c[15] ^ c[17] ^ c[19] ^ c[21] ^ c[22];
    newcrc[16] = d[255] ^ d[253] ^ d[251] ^ d[249] ^ d[247] ^ d[246] ^ d[243] ^ d[241] ^ d[240] ^ d[238] ^ d[232] ^ d[229] ^ d[228] ^ d[226] ^ d[225] ^ d[221] ^ d[220] ^ d[216] ^ d[214] ^ d[213] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[196] ^ d[194] ^ d[191] ^ d[189] ^ d[188] ^ d[186] ^ d[176] ^ d[175] ^ d[174] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[160] ^ d[159] ^ d[158] ^ d[157] ^ d[156] ^ d[155] ^ d[153] ^ d[152] ^ d[150] ^ d[143] ^ d[141] ^ d[139] ^ d[135] ^ d[134] ^ d[133] ^ d[131] ^ d[128] ^ d[126] ^ d[124] ^ d[120] ^ d[116] ^ d[112] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[102] ^ d[100] ^ d[95] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[81] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[70] ^ d[69] ^ d[68] ^ d[66] ^ d[64] ^ d[63] ^ d[60] ^ d[58] ^ d[55] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[45] ^ d[44] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[35] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[27] ^ d[25] ^ d[21] ^ d[20] ^ d[17] ^ d[13] ^ d[12] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[2] ^ c[5] ^ c[7] ^ c[8] ^ c[10] ^ c[13] ^ c[14] ^ c[16] ^ c[18] ^ c[20] ^ c[22];
    newcrc[17] = d[255] ^ d[250] ^ d[249] ^ d[247] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[238] ^ d[236] ^ d[235] ^ d[233] ^ d[232] ^ d[231] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[221] ^ d[219] ^ d[218] ^ d[214] ^ d[213] ^ d[211] ^ d[210] ^ d[207] ^ d[206] ^ d[204] ^ d[202] ^ d[201] ^ d[200] ^ d[197] ^ d[194] ^ d[193] ^ d[192] ^ d[187] ^ d[184] ^ d[178] ^ d[177] ^ d[175] ^ d[172] ^ d[171] ^ d[167] ^ d[166] ^ d[164] ^ d[162] ^ d[161] ^ d[160] ^ d[159] ^ d[157] ^ d[156] ^ d[153] ^ d[152] ^ d[151] ^ d[148] ^ d[147] ^ d[143] ^ d[139] ^ d[137] ^ d[135] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[128] ^ d[126] ^ d[124] ^ d[122] ^ d[119] ^ d[115] ^ d[114] ^ d[112] ^ d[110] ^ d[109] ^ d[105] ^ d[101] ^ d[98] ^ d[95] ^ d[94] ^ d[93] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[85] ^ d[83] ^ d[82] ^ d[81] ^ d[76] ^ d[75] ^ d[74] ^ d[72] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[64] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[45] ^ d[44] ^ d[42] ^ d[41] ^ d[40] ^ d[36] ^ d[33] ^ d[32] ^ d[30] ^ d[28] ^ d[23] ^ d[22] ^ d[15] ^ d[14] ^ d[8] ^ d[7] ^ d[5] ^ d[3] ^ d[0] ^ c[0] ^ c[2] ^ c[3] ^ c[5] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[22];
    newcrc[18] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[250] ^ d[249] ^ d[247] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[233] ^ d[231] ^ d[230] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[220] ^ d[218] ^ d[217] ^ d[214] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[206] ^ d[205] ^ d[202] ^ d[201] ^ d[198] ^ d[190] ^ d[189] ^ d[188] ^ d[185] ^ d[184] ^ d[179] ^ d[173] ^ d[171] ^ d[167] ^ d[166] ^ d[163] ^ d[161] ^ d[160] ^ d[157] ^ d[153] ^ d[149] ^ d[147] ^ d[143] ^ d[142] ^ d[139] ^ d[138] ^ d[137] ^ d[135] ^ d[134] ^ d[132] ^ d[131] ^ d[128] ^ d[126] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[117] ^ d[116] ^ d[114] ^ d[112] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[104] ^ d[103] ^ d[102] ^ d[99] ^ d[98] ^ d[93] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[87] ^ d[82] ^ d[81] ^ d[79] ^ d[78] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[63] ^ d[61] ^ d[60] ^ d[57] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[45] ^ d[44] ^ d[41] ^ d[39] ^ d[38] ^ d[37] ^ d[34] ^ d[33] ^ d[26] ^ d[24] ^ d[21] ^ d[18] ^ d[16] ^ d[13] ^ d[10] ^ d[8] ^ d[5] ^ d[4] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[14] ^ c[16] ^ c[17] ^ c[18] ^ c[19] ^ c[21] ^ c[22];
    newcrc[19] = d[255] ^ d[253] ^ d[252] ^ d[251] ^ d[250] ^ d[248] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[239] ^ d[238] ^ d[236] ^ d[235] ^ d[234] ^ d[232] ^ d[231] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[221] ^ d[219] ^ d[218] ^ d[215] ^ d[214] ^ d[213] ^ d[211] ^ d[209] ^ d[207] ^ d[206] ^ d[203] ^ d[202] ^ d[199] ^ d[191] ^ d[190] ^ d[189] ^ d[186] ^ d[185] ^ d[180] ^ d[174] ^ d[172] ^ d[168] ^ d[167] ^ d[164] ^ d[162] ^ d[161] ^ d[158] ^ d[154] ^ d[150] ^ d[148] ^ d[144] ^ d[143] ^ d[140] ^ d[139] ^ d[138] ^ d[136] ^ d[135] ^ d[133] ^ d[132] ^ d[129] ^ d[127] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[118] ^ d[117] ^ d[115] ^ d[113] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[103] ^ d[100] ^ d[99] ^ d[94] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[88] ^ d[83] ^ d[82] ^ d[80] ^ d[79] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[64] ^ d[62] ^ d[61] ^ d[58] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[46] ^ d[45] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[35] ^ d[34] ^ d[27] ^ d[25] ^ d[22] ^ d[19] ^ d[17] ^ d[14] ^ d[11] ^ d[9] ^ d[6] ^ d[5] ^ d[2] ^ d[1] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[15] ^ c[17] ^ c[18] ^ c[19] ^ c[20] ^ c[22];
    newcrc[20] = d[254] ^ d[253] ^ d[252] ^ d[251] ^ d[249] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[240] ^ d[239] ^ d[237] ^ d[236] ^ d[235] ^ d[233] ^ d[232] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[225] ^ d[222] ^ d[220] ^ d[219] ^ d[216] ^ d[215] ^ d[214] ^ d[212] ^ d[210] ^ d[208] ^ d[207] ^ d[204] ^ d[203] ^ d[200] ^ d[192] ^ d[191] ^ d[190] ^ d[187] ^ d[186] ^ d[181] ^ d[175] ^ d[173] ^ d[169] ^ d[168] ^ d[165] ^ d[163] ^ d[162] ^ d[159] ^ d[155] ^ d[151] ^ d[149] ^ d[145] ^ d[144] ^ d[141] ^ d[140] ^ d[139] ^ d[137] ^ d[136] ^ d[134] ^ d[133] ^ d[130] ^ d[128] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[119] ^ d[118] ^ d[116] ^ d[114] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[101] ^ d[100] ^ d[95] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[89] ^ d[84] ^ d[83] ^ d[81] ^ d[80] ^ d[78] ^ d[76] ^ d[75] ^ d[74] ^ d[72] ^ d[71] ^ d[69] ^ d[68] ^ d[65] ^ d[63] ^ d[62] ^ d[59] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[47] ^ d[46] ^ d[43] ^ d[41] ^ d[40] ^ d[39] ^ d[36] ^ d[35] ^ d[28] ^ d[26] ^ d[23] ^ d[20] ^ d[18] ^ d[15] ^ d[12] ^ d[10] ^ d[7] ^ d[6] ^ d[3] ^ d[2] ^ c[0] ^ c[2] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[12] ^ c[13] ^ c[16] ^ c[18] ^ c[19] ^ c[20] ^ c[21];
    newcrc[21] = d[255] ^ d[254] ^ d[253] ^ d[252] ^ d[250] ^ d[247] ^ d[246] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[238] ^ d[237] ^ d[236] ^ d[234] ^ d[233] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[226] ^ d[223] ^ d[221] ^ d[220] ^ d[217] ^ d[216] ^ d[215] ^ d[213] ^ d[211] ^ d[209] ^ d[208] ^ d[205] ^ d[204] ^ d[201] ^ d[193] ^ d[192] ^ d[191] ^ d[188] ^ d[187] ^ d[182] ^ d[176] ^ d[174] ^ d[170] ^ d[169] ^ d[166] ^ d[164] ^ d[163] ^ d[160] ^ d[156] ^ d[152] ^ d[150] ^ d[146] ^ d[145] ^ d[142] ^ d[141] ^ d[140] ^ d[138] ^ d[137] ^ d[135] ^ d[134] ^ d[131] ^ d[129] ^ d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[122] ^ d[120] ^ d[119] ^ d[117] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[102] ^ d[101] ^ d[96] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[90] ^ d[85] ^ d[84] ^ d[82] ^ d[81] ^ d[79] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[66] ^ d[64] ^ d[63] ^ d[60] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[48] ^ d[47] ^ d[44] ^ d[42] ^ d[41] ^ d[40] ^ d[37] ^ d[36] ^ d[29] ^ d[27] ^ d[24] ^ d[21] ^ d[19] ^ d[16] ^ d[13] ^ d[11] ^ d[8] ^ d[7] ^ d[4] ^ d[3] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[13] ^ c[14] ^ c[17] ^ c[19] ^ c[20] ^ c[21] ^ c[22];
    newcrc[22] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[248] ^ d[247] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[239] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[231] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[224] ^ d[222] ^ d[221] ^ d[218] ^ d[217] ^ d[216] ^ d[214] ^ d[212] ^ d[210] ^ d[209] ^ d[206] ^ d[205] ^ d[202] ^ d[194] ^ d[193] ^ d[192] ^ d[189] ^ d[188] ^ d[183] ^ d[177] ^ d[175] ^ d[171] ^ d[170] ^ d[167] ^ d[165] ^ d[164] ^ d[161] ^ d[157] ^ d[153] ^ d[151] ^ d[147] ^ d[146] ^ d[143] ^ d[142] ^ d[141] ^ d[139] ^ d[138] ^ d[136] ^ d[135] ^ d[132] ^ d[130] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[124] ^ d[123] ^ d[121] ^ d[120] ^ d[118] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[106] ^ d[103] ^ d[102] ^ d[97] ^ d[95] ^ d[94] ^ d[93] ^ d[92] ^ d[91] ^ d[86] ^ d[85] ^ d[83] ^ d[82] ^ d[80] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[71] ^ d[70] ^ d[67] ^ d[65] ^ d[64] ^ d[61] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[49] ^ d[48] ^ d[45] ^ d[43] ^ d[42] ^ d[41] ^ d[38] ^ d[37] ^ d[30] ^ d[28] ^ d[25] ^ d[22] ^ d[20] ^ d[17] ^ d[14] ^ d[12] ^ d[9] ^ d[8] ^ d[5] ^ d[4] ^ c[1] ^ c[2] ^ c[4] ^ c[5] ^ c[6] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[14] ^ c[15] ^ c[18] ^ c[20] ^ c[21] ^ c[22];
    crcf1 = newcrc;
  end
  endfunction


////////////////////////////////////////////////////////////////////////////////
// Copyright (C) 1999-2008 Easics NV.
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//
// Purpose : synthesizable CRC function
//   * polynomial: (0 1 3 6 7 8 10 11 13 14 16 18 19 20 22)
//   * data width: 256
//
// Info : tools@easics.be
//        http://www.easics.com
////////////////////////////////////////////////////////////////////////////////

  // polynomial: (0 1 3 6 7 8 10 11 13 14 16 18 19 20 22)
  // data width: 256
  // convention: the first serial bit is D[255]
  function [21:0] crcf0;

    input [255:0] Data;
    input [21:0] crc;
    reg [255:0] d;
    reg [21:0] c;
    reg [21:0] newcrc;
  begin
    d = Data;
    c = crc;

    newcrc[0] = d[255] ^ d[253] ^ d[252] ^ d[250] ^ d[249] ^ d[246] ^ d[245] ^ d[243] ^ d[242] ^ d[241] ^ d[239] ^ d[238] ^ d[237] ^ d[236] ^ d[233] ^ d[232] ^ d[228] ^ d[227] ^ d[226] ^ d[224] ^ d[222] ^ d[221] ^ d[220] ^ d[216] ^ d[215] ^ d[211] ^ d[208] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[195] ^ d[193] ^ d[192] ^ d[191] ^ d[190] ^ d[188] ^ d[182] ^ d[181] ^ d[179] ^ d[176] ^ d[175] ^ d[174] ^ d[172] ^ d[170] ^ d[165] ^ d[162] ^ d[160] ^ d[154] ^ d[150] ^ d[148] ^ d[147] ^ d[146] ^ d[145] ^ d[143] ^ d[138] ^ d[136] ^ d[135] ^ d[128] ^ d[127] ^ d[126] ^ d[124] ^ d[123] ^ d[122] ^ d[119] ^ d[116] ^ d[114] ^ d[112] ^ d[110] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[100] ^ d[99] ^ d[98] ^ d[87] ^ d[85] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[72] ^ d[71] ^ d[70] ^ d[66] ^ d[65] ^ d[63] ^ d[61] ^ d[59] ^ d[58] ^ d[56] ^ d[55] ^ d[54] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[47] ^ d[45] ^ d[44] ^ d[43] ^ d[42] ^ d[40] ^ d[39] ^ d[37] ^ d[33] ^ d[32] ^ d[31] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[16] ^ d[13] ^ d[11] ^ d[8] ^ d[7] ^ d[6] ^ d[3] ^ d[2] ^ d[0] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[15] ^ c[16] ^ c[18] ^ c[19] ^ c[21];
    newcrc[1] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[249] ^ d[247] ^ d[245] ^ d[244] ^ d[241] ^ d[240] ^ d[236] ^ d[234] ^ d[232] ^ d[229] ^ d[226] ^ d[225] ^ d[224] ^ d[223] ^ d[220] ^ d[217] ^ d[215] ^ d[212] ^ d[211] ^ d[209] ^ d[208] ^ d[206] ^ d[199] ^ d[196] ^ d[195] ^ d[194] ^ d[190] ^ d[189] ^ d[188] ^ d[183] ^ d[181] ^ d[180] ^ d[179] ^ d[177] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[170] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[161] ^ d[160] ^ d[155] ^ d[154] ^ d[151] ^ d[150] ^ d[149] ^ d[145] ^ d[144] ^ d[143] ^ d[139] ^ d[138] ^ d[137] ^ d[135] ^ d[129] ^ d[126] ^ d[125] ^ d[122] ^ d[120] ^ d[119] ^ d[117] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[110] ^ d[108] ^ d[104] ^ d[101] ^ d[98] ^ d[88] ^ d[87] ^ d[86] ^ d[85] ^ d[82] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[70] ^ d[67] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[53] ^ d[52] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[42] ^ d[41] ^ d[39] ^ d[38] ^ d[37] ^ d[34] ^ d[31] ^ d[28] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[12] ^ d[11] ^ d[9] ^ d[6] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[2] ^ c[6] ^ c[7] ^ c[10] ^ c[11] ^ c[13] ^ c[15] ^ c[17] ^ c[18] ^ c[20] ^ c[21];
    newcrc[2] = d[255] ^ d[253] ^ d[252] ^ d[250] ^ d[248] ^ d[246] ^ d[245] ^ d[242] ^ d[241] ^ d[237] ^ d[235] ^ d[233] ^ d[230] ^ d[227] ^ d[226] ^ d[225] ^ d[224] ^ d[221] ^ d[218] ^ d[216] ^ d[213] ^ d[212] ^ d[210] ^ d[209] ^ d[207] ^ d[200] ^ d[197] ^ d[196] ^ d[195] ^ d[191] ^ d[190] ^ d[189] ^ d[184] ^ d[182] ^ d[181] ^ d[180] ^ d[178] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[156] ^ d[155] ^ d[152] ^ d[151] ^ d[150] ^ d[146] ^ d[145] ^ d[144] ^ d[140] ^ d[139] ^ d[138] ^ d[136] ^ d[130] ^ d[127] ^ d[126] ^ d[123] ^ d[121] ^ d[120] ^ d[118] ^ d[117] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[111] ^ d[109] ^ d[105] ^ d[102] ^ d[99] ^ d[89] ^ d[88] ^ d[87] ^ d[86] ^ d[83] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[71] ^ d[68] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[59] ^ d[58] ^ d[54] ^ d[53] ^ d[50] ^ d[49] ^ d[48] ^ d[47] ^ d[43] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[35] ^ d[32] ^ d[29] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[14] ^ d[13] ^ d[12] ^ d[10] ^ d[7] ^ d[5] ^ d[3] ^ d[2] ^ d[1] ^ c[1] ^ c[3] ^ c[7] ^ c[8] ^ c[11] ^ c[12] ^ c[14] ^ c[16] ^ c[18] ^ c[19] ^ c[21];
    newcrc[3] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[250] ^ d[247] ^ d[245] ^ d[241] ^ d[239] ^ d[237] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[225] ^ d[224] ^ d[221] ^ d[220] ^ d[219] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[213] ^ d[210] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[195] ^ d[193] ^ d[188] ^ d[185] ^ d[183] ^ d[173] ^ d[170] ^ d[168] ^ d[167] ^ d[164] ^ d[163] ^ d[160] ^ d[157] ^ d[156] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[150] ^ d[148] ^ d[143] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[135] ^ d[131] ^ d[126] ^ d[123] ^ d[121] ^ d[118] ^ d[117] ^ d[115] ^ d[113] ^ d[107] ^ d[105] ^ d[104] ^ d[103] ^ d[99] ^ d[98] ^ d[90] ^ d[89] ^ d[88] ^ d[85] ^ d[84] ^ d[81] ^ d[80] ^ d[71] ^ d[70] ^ d[69] ^ d[67] ^ d[64] ^ d[62] ^ d[61] ^ d[60] ^ d[58] ^ d[56] ^ d[53] ^ d[48] ^ d[47] ^ d[45] ^ d[42] ^ d[41] ^ d[37] ^ d[36] ^ d[32] ^ d[31] ^ d[30] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[15] ^ d[14] ^ d[7] ^ d[4] ^ d[0] ^ c[0] ^ c[3] ^ c[5] ^ c[7] ^ c[11] ^ c[13] ^ c[16] ^ c[17] ^ c[18] ^ c[20] ^ c[21];
    newcrc[4] = d[255] ^ d[253] ^ d[252] ^ d[251] ^ d[248] ^ d[246] ^ d[242] ^ d[240] ^ d[238] ^ d[235] ^ d[234] ^ d[233] ^ d[232] ^ d[226] ^ d[225] ^ d[222] ^ d[221] ^ d[220] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[214] ^ d[211] ^ d[206] ^ d[205] ^ d[204] ^ d[203] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[194] ^ d[189] ^ d[186] ^ d[184] ^ d[174] ^ d[171] ^ d[169] ^ d[168] ^ d[165] ^ d[164] ^ d[161] ^ d[158] ^ d[157] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[149] ^ d[144] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[136] ^ d[132] ^ d[127] ^ d[124] ^ d[122] ^ d[119] ^ d[118] ^ d[116] ^ d[114] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[100] ^ d[99] ^ d[91] ^ d[90] ^ d[89] ^ d[86] ^ d[85] ^ d[82] ^ d[81] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[65] ^ d[63] ^ d[62] ^ d[61] ^ d[59] ^ d[57] ^ d[54] ^ d[49] ^ d[48] ^ d[46] ^ d[43] ^ d[42] ^ d[38] ^ d[37] ^ d[33] ^ d[32] ^ d[31] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[16] ^ d[15] ^ d[8] ^ d[5] ^ d[1] ^ c[0] ^ c[1] ^ c[4] ^ c[6] ^ c[8] ^ c[12] ^ c[14] ^ c[17] ^ c[18] ^ c[19] ^ c[21];
    newcrc[5] = d[254] ^ d[253] ^ d[252] ^ d[249] ^ d[247] ^ d[243] ^ d[241] ^ d[239] ^ d[236] ^ d[235] ^ d[234] ^ d[233] ^ d[227] ^ d[226] ^ d[223] ^ d[222] ^ d[221] ^ d[219] ^ d[218] ^ d[217] ^ d[216] ^ d[215] ^ d[212] ^ d[207] ^ d[206] ^ d[205] ^ d[204] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[195] ^ d[190] ^ d[187] ^ d[185] ^ d[175] ^ d[172] ^ d[170] ^ d[169] ^ d[166] ^ d[165] ^ d[162] ^ d[159] ^ d[158] ^ d[156] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[150] ^ d[145] ^ d[143] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[138] ^ d[137] ^ d[133] ^ d[128] ^ d[125] ^ d[123] ^ d[120] ^ d[119] ^ d[117] ^ d[115] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[101] ^ d[100] ^ d[92] ^ d[91] ^ d[90] ^ d[87] ^ d[86] ^ d[83] ^ d[82] ^ d[73] ^ d[72] ^ d[71] ^ d[69] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[60] ^ d[58] ^ d[55] ^ d[50] ^ d[49] ^ d[47] ^ d[44] ^ d[43] ^ d[39] ^ d[38] ^ d[34] ^ d[33] ^ d[32] ^ d[29] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[17] ^ d[16] ^ d[9] ^ d[6] ^ d[2] ^ c[0] ^ c[1] ^ c[2] ^ c[5] ^ c[7] ^ c[9] ^ c[13] ^ c[15] ^ c[18] ^ c[19] ^ c[20];
    newcrc[6] = d[254] ^ d[252] ^ d[249] ^ d[248] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[235] ^ d[234] ^ d[233] ^ d[232] ^ d[226] ^ d[223] ^ d[221] ^ d[219] ^ d[218] ^ d[217] ^ d[215] ^ d[213] ^ d[211] ^ d[207] ^ d[206] ^ d[204] ^ d[198] ^ d[196] ^ d[195] ^ d[193] ^ d[192] ^ d[190] ^ d[186] ^ d[182] ^ d[181] ^ d[179] ^ d[175] ^ d[174] ^ d[173] ^ d[172] ^ d[171] ^ d[167] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[159] ^ d[157] ^ d[156] ^ d[155] ^ d[153] ^ d[151] ^ d[150] ^ d[148] ^ d[147] ^ d[145] ^ d[144] ^ d[142] ^ d[141] ^ d[140] ^ d[139] ^ d[136] ^ d[135] ^ d[134] ^ d[129] ^ d[128] ^ d[127] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[119] ^ d[118] ^ d[114] ^ d[112] ^ d[108] ^ d[105] ^ d[104] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[93] ^ d[92] ^ d[91] ^ d[88] ^ d[85] ^ d[84] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[71] ^ d[67] ^ d[66] ^ d[64] ^ d[58] ^ d[55] ^ d[54] ^ d[53] ^ d[49] ^ d[48] ^ d[47] ^ d[43] ^ d[42] ^ d[37] ^ d[35] ^ d[34] ^ d[32] ^ d[31] ^ d[30] ^ d[29] ^ d[28] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[17] ^ d[16] ^ d[13] ^ d[11] ^ d[10] ^ d[8] ^ d[6] ^ d[2] ^ d[0] ^ c[0] ^ c[1] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[14] ^ c[15] ^ c[18] ^ c[20];
    newcrc[7] = d[252] ^ d[247] ^ d[244] ^ d[243] ^ d[240] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[232] ^ d[228] ^ d[226] ^ d[221] ^ d[219] ^ d[218] ^ d[215] ^ d[214] ^ d[212] ^ d[211] ^ d[207] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[197] ^ d[196] ^ d[195] ^ d[194] ^ d[192] ^ d[190] ^ d[188] ^ d[187] ^ d[183] ^ d[181] ^ d[180] ^ d[179] ^ d[173] ^ d[170] ^ d[168] ^ d[167] ^ d[166] ^ d[165] ^ d[164] ^ d[163] ^ d[162] ^ d[158] ^ d[157] ^ d[156] ^ d[152] ^ d[151] ^ d[150] ^ d[149] ^ d[147] ^ d[142] ^ d[141] ^ d[140] ^ d[138] ^ d[137] ^ d[130] ^ d[129] ^ d[127] ^ d[126] ^ d[121] ^ d[120] ^ d[116] ^ d[115] ^ d[114] ^ d[113] ^ d[112] ^ d[110] ^ d[109] ^ d[107] ^ d[104] ^ d[103] ^ d[102] ^ d[101] ^ d[98] ^ d[94] ^ d[93] ^ d[92] ^ d[89] ^ d[87] ^ d[86] ^ d[84] ^ d[82] ^ d[77] ^ d[76] ^ d[74] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[66] ^ d[63] ^ d[61] ^ d[58] ^ d[53] ^ d[51] ^ d[48] ^ d[47] ^ d[45] ^ d[42] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[30] ^ d[29] ^ d[27] ^ d[26] ^ d[25] ^ d[19] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[12] ^ d[9] ^ d[8] ^ d[6] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[6] ^ c[9] ^ c[10] ^ c[13] ^ c[18];
    newcrc[8] = d[255] ^ d[252] ^ d[250] ^ d[249] ^ d[248] ^ d[246] ^ d[244] ^ d[243] ^ d[242] ^ d[237] ^ d[235] ^ d[232] ^ d[229] ^ d[228] ^ d[226] ^ d[224] ^ d[221] ^ d[219] ^ d[213] ^ d[212] ^ d[211] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[196] ^ d[192] ^ d[190] ^ d[189] ^ d[184] ^ d[180] ^ d[179] ^ d[176] ^ d[175] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[162] ^ d[160] ^ d[159] ^ d[158] ^ d[157] ^ d[154] ^ d[153] ^ d[152] ^ d[151] ^ d[147] ^ d[146] ^ d[145] ^ d[142] ^ d[141] ^ d[139] ^ d[136] ^ d[135] ^ d[131] ^ d[130] ^ d[126] ^ d[124] ^ d[123] ^ d[121] ^ d[119] ^ d[117] ^ d[115] ^ d[113] ^ d[112] ^ d[111] ^ d[108] ^ d[107] ^ d[106] ^ d[103] ^ d[102] ^ d[100] ^ d[98] ^ d[95] ^ d[94] ^ d[93] ^ d[90] ^ d[88] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[58] ^ d[56] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[44] ^ d[42] ^ d[41] ^ d[38] ^ d[36] ^ d[33] ^ d[32] ^ d[30] ^ d[28] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[19] ^ d[17] ^ d[16] ^ d[15] ^ d[14] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[6] ^ d[1] ^ d[0] ^ c[1] ^ c[3] ^ c[8] ^ c[9] ^ c[10] ^ c[12] ^ c[14] ^ c[15] ^ c[16] ^ c[18] ^ c[21];
    newcrc[9] = d[253] ^ d[251] ^ d[250] ^ d[249] ^ d[247] ^ d[245] ^ d[244] ^ d[243] ^ d[238] ^ d[236] ^ d[233] ^ d[230] ^ d[229] ^ d[227] ^ d[225] ^ d[222] ^ d[220] ^ d[214] ^ d[213] ^ d[212] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[193] ^ d[191] ^ d[190] ^ d[185] ^ d[181] ^ d[180] ^ d[177] ^ d[176] ^ d[173] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[168] ^ d[167] ^ d[165] ^ d[164] ^ d[163] ^ d[161] ^ d[160] ^ d[159] ^ d[158] ^ d[155] ^ d[154] ^ d[153] ^ d[152] ^ d[148] ^ d[147] ^ d[146] ^ d[143] ^ d[142] ^ d[140] ^ d[137] ^ d[136] ^ d[132] ^ d[131] ^ d[127] ^ d[125] ^ d[124] ^ d[122] ^ d[120] ^ d[118] ^ d[116] ^ d[114] ^ d[113] ^ d[112] ^ d[109] ^ d[108] ^ d[107] ^ d[104] ^ d[103] ^ d[101] ^ d[99] ^ d[96] ^ d[95] ^ d[94] ^ d[91] ^ d[89] ^ d[84] ^ d[82] ^ d[81] ^ d[80] ^ d[71] ^ d[70] ^ d[69] ^ d[68] ^ d[67] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[59] ^ d[57] ^ d[56] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[39] ^ d[37] ^ d[34] ^ d[33] ^ d[31] ^ d[29] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[20] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[7] ^ d[2] ^ d[1] ^ c[2] ^ c[4] ^ c[9] ^ c[10] ^ c[11] ^ c[13] ^ c[15] ^ c[16] ^ c[17] ^ c[19];
    newcrc[10] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[249] ^ d[248] ^ d[244] ^ d[243] ^ d[242] ^ d[241] ^ d[238] ^ d[236] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[227] ^ d[224] ^ d[223] ^ d[222] ^ d[220] ^ d[216] ^ d[214] ^ d[213] ^ d[211] ^ d[208] ^ d[205] ^ d[204] ^ d[203] ^ d[198] ^ d[195] ^ d[194] ^ d[193] ^ d[190] ^ d[188] ^ d[186] ^ d[179] ^ d[178] ^ d[177] ^ d[176] ^ d[175] ^ d[173] ^ d[171] ^ d[169] ^ d[168] ^ d[166] ^ d[164] ^ d[161] ^ d[159] ^ d[156] ^ d[155] ^ d[153] ^ d[150] ^ d[149] ^ d[146] ^ d[145] ^ d[144] ^ d[141] ^ d[137] ^ d[136] ^ d[135] ^ d[133] ^ d[132] ^ d[127] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[117] ^ d[116] ^ d[115] ^ d[113] ^ d[112] ^ d[109] ^ d[108] ^ d[107] ^ d[106] ^ d[102] ^ d[99] ^ d[98] ^ d[97] ^ d[96] ^ d[95] ^ d[92] ^ d[90] ^ d[87] ^ d[83] ^ d[82] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[69] ^ d[68] ^ d[67] ^ d[64] ^ d[61] ^ d[60] ^ d[59] ^ d[57] ^ d[56] ^ d[52] ^ d[51] ^ d[48] ^ d[46] ^ d[45] ^ d[42] ^ d[39] ^ d[38] ^ d[37] ^ d[35] ^ d[34] ^ d[33] ^ d[31] ^ d[30] ^ d[22] ^ d[20] ^ d[17] ^ d[12] ^ d[10] ^ d[7] ^ d[6] ^ d[0] ^ c[0] ^ c[2] ^ c[4] ^ c[7] ^ c[8] ^ c[9] ^ c[10] ^ c[14] ^ c[15] ^ c[17] ^ c[19] ^ c[20] ^ c[21];
    newcrc[11] = d[254] ^ d[253] ^ d[246] ^ d[244] ^ d[241] ^ d[238] ^ d[236] ^ d[235] ^ d[234] ^ d[231] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[222] ^ d[220] ^ d[217] ^ d[216] ^ d[214] ^ d[212] ^ d[211] ^ d[209] ^ d[208] ^ d[206] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[196] ^ d[194] ^ d[193] ^ d[192] ^ d[190] ^ d[189] ^ d[188] ^ d[187] ^ d[182] ^ d[181] ^ d[180] ^ d[178] ^ d[177] ^ d[175] ^ d[169] ^ d[167] ^ d[157] ^ d[156] ^ d[151] ^ d[148] ^ d[143] ^ d[142] ^ d[137] ^ d[135] ^ d[134] ^ d[133] ^ d[127] ^ d[125] ^ d[124] ^ d[119] ^ d[118] ^ d[117] ^ d[113] ^ d[112] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[97] ^ d[96] ^ d[93] ^ d[91] ^ d[88] ^ d[87] ^ d[85] ^ d[84] ^ d[83] ^ d[77] ^ d[76] ^ d[75] ^ d[72] ^ d[71] ^ d[69] ^ d[68] ^ d[66] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[57] ^ d[56] ^ d[55] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[46] ^ d[45] ^ d[44] ^ d[42] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[27] ^ d[26] ^ d[25] ^ d[24] ^ d[22] ^ d[20] ^ d[19] ^ d[16] ^ d[6] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[4] ^ c[7] ^ c[10] ^ c[12] ^ c[19] ^ c[20];
    newcrc[12] = d[255] ^ d[254] ^ d[247] ^ d[245] ^ d[242] ^ d[239] ^ d[237] ^ d[236] ^ d[235] ^ d[232] ^ d[228] ^ d[227] ^ d[226] ^ d[224] ^ d[223] ^ d[221] ^ d[218] ^ d[217] ^ d[215] ^ d[213] ^ d[212] ^ d[210] ^ d[209] ^ d[207] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[197] ^ d[195] ^ d[194] ^ d[193] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[183] ^ d[182] ^ d[181] ^ d[179] ^ d[178] ^ d[176] ^ d[170] ^ d[168] ^ d[158] ^ d[157] ^ d[152] ^ d[149] ^ d[144] ^ d[143] ^ d[138] ^ d[136] ^ d[135] ^ d[134] ^ d[128] ^ d[126] ^ d[125] ^ d[120] ^ d[119] ^ d[118] ^ d[114] ^ d[113] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[105] ^ d[104] ^ d[98] ^ d[97] ^ d[94] ^ d[92] ^ d[89] ^ d[88] ^ d[86] ^ d[85] ^ d[84] ^ d[78] ^ d[77] ^ d[76] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[67] ^ d[64] ^ d[63] ^ d[61] ^ d[60] ^ d[58] ^ d[57] ^ d[56] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[23] ^ d[21] ^ d[20] ^ d[17] ^ d[7] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[8] ^ c[11] ^ c[13] ^ c[20] ^ c[21];
    newcrc[13] = d[253] ^ d[252] ^ d[250] ^ d[249] ^ d[248] ^ d[245] ^ d[242] ^ d[241] ^ d[240] ^ d[239] ^ d[232] ^ d[229] ^ d[226] ^ d[225] ^ d[221] ^ d[220] ^ d[219] ^ d[218] ^ d[215] ^ d[214] ^ d[213] ^ d[210] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[196] ^ d[194] ^ d[193] ^ d[189] ^ d[188] ^ d[184] ^ d[183] ^ d[181] ^ d[180] ^ d[177] ^ d[176] ^ d[175] ^ d[174] ^ d[172] ^ d[171] ^ d[170] ^ d[169] ^ d[165] ^ d[162] ^ d[160] ^ d[159] ^ d[158] ^ d[154] ^ d[153] ^ d[148] ^ d[147] ^ d[146] ^ d[144] ^ d[143] ^ d[139] ^ d[138] ^ d[137] ^ d[129] ^ d[128] ^ d[124] ^ d[123] ^ d[122] ^ d[121] ^ d[120] ^ d[116] ^ d[115] ^ d[112] ^ d[111] ^ d[108] ^ d[104] ^ d[100] ^ d[95] ^ d[93] ^ d[90] ^ d[89] ^ d[86] ^ d[81] ^ d[80] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[68] ^ d[66] ^ d[64] ^ d[63] ^ d[62] ^ d[57] ^ d[55] ^ d[52] ^ d[51] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[45] ^ d[43] ^ d[42] ^ d[38] ^ d[36] ^ d[35] ^ d[33] ^ d[32] ^ d[31] ^ d[29] ^ d[28] ^ d[25] ^ d[23] ^ d[20] ^ d[19] ^ d[16] ^ d[13] ^ d[11] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[0] ^ c[5] ^ c[6] ^ c[7] ^ c[8] ^ c[11] ^ c[14] ^ c[15] ^ c[16] ^ c[18] ^ c[19];
    newcrc[14] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[245] ^ d[240] ^ d[239] ^ d[238] ^ d[237] ^ d[236] ^ d[232] ^ d[230] ^ d[228] ^ d[224] ^ d[219] ^ d[214] ^ d[208] ^ d[205] ^ d[204] ^ d[203] ^ d[197] ^ d[194] ^ d[193] ^ d[192] ^ d[191] ^ d[189] ^ d[188] ^ d[185] ^ d[184] ^ d[179] ^ d[178] ^ d[177] ^ d[174] ^ d[173] ^ d[171] ^ d[166] ^ d[165] ^ d[163] ^ d[162] ^ d[161] ^ d[159] ^ d[155] ^ d[150] ^ d[149] ^ d[146] ^ d[144] ^ d[143] ^ d[140] ^ d[139] ^ d[136] ^ d[135] ^ d[130] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[125] ^ d[121] ^ d[119] ^ d[117] ^ d[114] ^ d[113] ^ d[110] ^ d[109] ^ d[107] ^ d[106] ^ d[104] ^ d[101] ^ d[100] ^ d[99] ^ d[98] ^ d[96] ^ d[94] ^ d[91] ^ d[90] ^ d[85] ^ d[82] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[64] ^ d[61] ^ d[59] ^ d[55] ^ d[54] ^ d[52] ^ d[46] ^ d[45] ^ d[42] ^ d[40] ^ d[36] ^ d[34] ^ d[31] ^ d[30] ^ d[29] ^ d[27] ^ d[25] ^ d[23] ^ d[22] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[13] ^ d[12] ^ d[11] ^ d[5] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[2] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[11] ^ c[17] ^ c[18] ^ c[20] ^ c[21];
    newcrc[15] = d[255] ^ d[253] ^ d[252] ^ d[246] ^ d[241] ^ d[240] ^ d[239] ^ d[238] ^ d[237] ^ d[233] ^ d[231] ^ d[229] ^ d[225] ^ d[220] ^ d[215] ^ d[209] ^ d[206] ^ d[205] ^ d[204] ^ d[198] ^ d[195] ^ d[194] ^ d[193] ^ d[192] ^ d[190] ^ d[189] ^ d[186] ^ d[185] ^ d[180] ^ d[179] ^ d[178] ^ d[175] ^ d[174] ^ d[172] ^ d[167] ^ d[166] ^ d[164] ^ d[163] ^ d[162] ^ d[160] ^ d[156] ^ d[151] ^ d[150] ^ d[147] ^ d[145] ^ d[144] ^ d[141] ^ d[140] ^ d[137] ^ d[136] ^ d[131] ^ d[130] ^ d[129] ^ d[128] ^ d[127] ^ d[126] ^ d[122] ^ d[120] ^ d[118] ^ d[115] ^ d[114] ^ d[111] ^ d[110] ^ d[108] ^ d[107] ^ d[105] ^ d[102] ^ d[101] ^ d[100] ^ d[99] ^ d[97] ^ d[95] ^ d[92] ^ d[91] ^ d[86] ^ d[83] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[65] ^ d[62] ^ d[60] ^ d[56] ^ d[55] ^ d[53] ^ d[47] ^ d[46] ^ d[43] ^ d[41] ^ d[37] ^ d[35] ^ d[32] ^ d[31] ^ d[30] ^ d[28] ^ d[26] ^ d[24] ^ d[23] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[14] ^ d[13] ^ d[12] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ c[3] ^ c[4] ^ c[5] ^ c[6] ^ c[7] ^ c[12] ^ c[18] ^ c[19] ^ c[21];
    newcrc[16] = d[255] ^ d[254] ^ d[252] ^ d[250] ^ d[249] ^ d[247] ^ d[246] ^ d[245] ^ d[243] ^ d[240] ^ d[237] ^ d[236] ^ d[234] ^ d[233] ^ d[230] ^ d[228] ^ d[227] ^ d[224] ^ d[222] ^ d[220] ^ d[215] ^ d[211] ^ d[210] ^ d[208] ^ d[207] ^ d[206] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[196] ^ d[194] ^ d[192] ^ d[188] ^ d[187] ^ d[186] ^ d[182] ^ d[180] ^ d[174] ^ d[173] ^ d[172] ^ d[170] ^ d[168] ^ d[167] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[160] ^ d[157] ^ d[154] ^ d[152] ^ d[151] ^ d[150] ^ d[147] ^ d[143] ^ d[142] ^ d[141] ^ d[137] ^ d[136] ^ d[135] ^ d[132] ^ d[131] ^ d[130] ^ d[129] ^ d[126] ^ d[124] ^ d[122] ^ d[121] ^ d[115] ^ d[114] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[107] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[101] ^ d[99] ^ d[96] ^ d[93] ^ d[92] ^ d[85] ^ d[84] ^ d[82] ^ d[77] ^ d[76] ^ d[74] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[65] ^ d[59] ^ d[58] ^ d[57] ^ d[55] ^ d[53] ^ d[51] ^ d[50] ^ d[49] ^ d[48] ^ d[45] ^ d[43] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[36] ^ d[29] ^ d[26] ^ d[23] ^ d[22] ^ d[15] ^ d[14] ^ d[11] ^ d[8] ^ d[6] ^ d[5] ^ d[4] ^ d[0] ^ c[0] ^ c[2] ^ c[3] ^ c[6] ^ c[9] ^ c[11] ^ c[12] ^ c[13] ^ c[15] ^ c[16] ^ c[18] ^ c[20] ^ c[21];
    newcrc[17] = d[255] ^ d[253] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[244] ^ d[241] ^ d[238] ^ d[237] ^ d[235] ^ d[234] ^ d[231] ^ d[229] ^ d[228] ^ d[225] ^ d[223] ^ d[221] ^ d[216] ^ d[212] ^ d[211] ^ d[209] ^ d[208] ^ d[207] ^ d[205] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[197] ^ d[195] ^ d[193] ^ d[189] ^ d[188] ^ d[187] ^ d[183] ^ d[181] ^ d[175] ^ d[174] ^ d[173] ^ d[171] ^ d[169] ^ d[168] ^ d[165] ^ d[164] ^ d[163] ^ d[162] ^ d[161] ^ d[158] ^ d[155] ^ d[153] ^ d[152] ^ d[151] ^ d[148] ^ d[144] ^ d[143] ^ d[142] ^ d[138] ^ d[137] ^ d[136] ^ d[133] ^ d[132] ^ d[131] ^ d[130] ^ d[127] ^ d[125] ^ d[123] ^ d[122] ^ d[116] ^ d[115] ^ d[112] ^ d[111] ^ d[110] ^ d[109] ^ d[108] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[100] ^ d[97] ^ d[94] ^ d[93] ^ d[86] ^ d[85] ^ d[83] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[66] ^ d[60] ^ d[59] ^ d[58] ^ d[56] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[49] ^ d[46] ^ d[44] ^ d[41] ^ d[40] ^ d[39] ^ d[38] ^ d[37] ^ d[30] ^ d[27] ^ d[24] ^ d[23] ^ d[16] ^ d[15] ^ d[12] ^ d[9] ^ d[7] ^ d[6] ^ d[5] ^ d[1] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[7] ^ c[10] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[21];
    newcrc[18] = d[255] ^ d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[243] ^ d[241] ^ d[237] ^ d[235] ^ d[233] ^ d[230] ^ d[229] ^ d[228] ^ d[227] ^ d[221] ^ d[220] ^ d[217] ^ d[216] ^ d[215] ^ d[213] ^ d[212] ^ d[211] ^ d[210] ^ d[209] ^ d[206] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[196] ^ d[195] ^ d[194] ^ d[193] ^ d[192] ^ d[191] ^ d[189] ^ d[184] ^ d[181] ^ d[179] ^ d[169] ^ d[166] ^ d[164] ^ d[163] ^ d[160] ^ d[159] ^ d[156] ^ d[153] ^ d[152] ^ d[150] ^ d[149] ^ d[148] ^ d[147] ^ d[146] ^ d[144] ^ d[139] ^ d[137] ^ d[136] ^ d[135] ^ d[134] ^ d[133] ^ d[132] ^ d[131] ^ d[127] ^ d[122] ^ d[119] ^ d[117] ^ d[114] ^ d[113] ^ d[111] ^ d[109] ^ d[103] ^ d[101] ^ d[100] ^ d[99] ^ d[95] ^ d[94] ^ d[86] ^ d[85] ^ d[84] ^ d[81] ^ d[80] ^ d[77] ^ d[76] ^ d[67] ^ d[66] ^ d[65] ^ d[63] ^ d[60] ^ d[58] ^ d[57] ^ d[56] ^ d[54] ^ d[52] ^ d[49] ^ d[44] ^ d[43] ^ d[41] ^ d[38] ^ d[37] ^ d[33] ^ d[32] ^ d[28] ^ d[27] ^ d[26] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[11] ^ d[10] ^ d[3] ^ d[0] ^ c[1] ^ c[3] ^ c[7] ^ c[9] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[20] ^ c[21];
    newcrc[19] = d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[246] ^ d[245] ^ d[244] ^ d[243] ^ d[241] ^ d[239] ^ d[237] ^ d[234] ^ d[233] ^ d[232] ^ d[231] ^ d[230] ^ d[229] ^ d[227] ^ d[226] ^ d[224] ^ d[220] ^ d[218] ^ d[217] ^ d[215] ^ d[214] ^ d[213] ^ d[212] ^ d[210] ^ d[208] ^ d[207] ^ d[205] ^ d[204] ^ d[203] ^ d[197] ^ d[196] ^ d[194] ^ d[191] ^ d[188] ^ d[185] ^ d[181] ^ d[180] ^ d[179] ^ d[176] ^ d[175] ^ d[174] ^ d[172] ^ d[167] ^ d[164] ^ d[162] ^ d[161] ^ d[157] ^ d[153] ^ d[151] ^ d[149] ^ d[146] ^ d[143] ^ d[140] ^ d[137] ^ d[134] ^ d[133] ^ d[132] ^ d[127] ^ d[126] ^ d[124] ^ d[122] ^ d[120] ^ d[119] ^ d[118] ^ d[116] ^ d[115] ^ d[107] ^ d[106] ^ d[105] ^ d[102] ^ d[101] ^ d[99] ^ d[98] ^ d[96] ^ d[95] ^ d[86] ^ d[82] ^ d[80] ^ d[79] ^ d[75] ^ d[72] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[65] ^ d[64] ^ d[63] ^ d[57] ^ d[56] ^ d[54] ^ d[51] ^ d[49] ^ d[47] ^ d[43] ^ d[40] ^ d[38] ^ d[37] ^ d[34] ^ d[32] ^ d[31] ^ d[29] ^ d[28] ^ d[26] ^ d[25] ^ d[16] ^ d[13] ^ d[12] ^ d[8] ^ d[7] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[0] ^ c[3] ^ c[5] ^ c[7] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[20];
    newcrc[20] = d[254] ^ d[253] ^ d[251] ^ d[250] ^ d[248] ^ d[247] ^ d[244] ^ d[243] ^ d[241] ^ d[240] ^ d[239] ^ d[237] ^ d[236] ^ d[235] ^ d[234] ^ d[231] ^ d[230] ^ d[226] ^ d[225] ^ d[224] ^ d[222] ^ d[220] ^ d[219] ^ d[218] ^ d[214] ^ d[213] ^ d[209] ^ d[206] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[197] ^ d[193] ^ d[191] ^ d[190] ^ d[189] ^ d[188] ^ d[186] ^ d[180] ^ d[179] ^ d[177] ^ d[174] ^ d[173] ^ d[172] ^ d[170] ^ d[168] ^ d[163] ^ d[160] ^ d[158] ^ d[152] ^ d[148] ^ d[146] ^ d[145] ^ d[144] ^ d[143] ^ d[141] ^ d[136] ^ d[134] ^ d[133] ^ d[126] ^ d[125] ^ d[124] ^ d[122] ^ d[121] ^ d[120] ^ d[117] ^ d[114] ^ d[112] ^ d[110] ^ d[108] ^ d[105] ^ d[104] ^ d[103] ^ d[102] ^ d[98] ^ d[97] ^ d[96] ^ d[85] ^ d[83] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[70] ^ d[69] ^ d[68] ^ d[64] ^ d[63] ^ d[61] ^ d[59] ^ d[57] ^ d[56] ^ d[54] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[45] ^ d[43] ^ d[42] ^ d[41] ^ d[40] ^ d[38] ^ d[37] ^ d[35] ^ d[31] ^ d[30] ^ d[29] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[14] ^ d[11] ^ d[9] ^ d[6] ^ d[5] ^ d[4] ^ d[1] ^ d[0] ^ c[0] ^ c[1] ^ c[2] ^ c[3] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[13] ^ c[14] ^ c[16] ^ c[17] ^ c[19] ^ c[20];
    newcrc[21] = d[255] ^ d[254] ^ d[252] ^ d[251] ^ d[249] ^ d[248] ^ d[245] ^ d[244] ^ d[242] ^ d[241] ^ d[240] ^ d[238] ^ d[237] ^ d[236] ^ d[235] ^ d[232] ^ d[231] ^ d[227] ^ d[226] ^ d[225] ^ d[223] ^ d[221] ^ d[220] ^ d[219] ^ d[215] ^ d[214] ^ d[210] ^ d[207] ^ d[204] ^ d[203] ^ d[202] ^ d[201] ^ d[200] ^ d[199] ^ d[198] ^ d[194] ^ d[192] ^ d[191] ^ d[190] ^ d[189] ^ d[187] ^ d[181] ^ d[180] ^ d[178] ^ d[175] ^ d[174] ^ d[173] ^ d[171] ^ d[169] ^ d[164] ^ d[161] ^ d[159] ^ d[153] ^ d[149] ^ d[147] ^ d[146] ^ d[145] ^ d[144] ^ d[142] ^ d[137] ^ d[135] ^ d[134] ^ d[127] ^ d[126] ^ d[125] ^ d[123] ^ d[122] ^ d[121] ^ d[118] ^ d[115] ^ d[113] ^ d[111] ^ d[109] ^ d[106] ^ d[105] ^ d[104] ^ d[103] ^ d[99] ^ d[98] ^ d[97] ^ d[86] ^ d[84] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[71] ^ d[70] ^ d[69] ^ d[65] ^ d[64] ^ d[62] ^ d[60] ^ d[58] ^ d[57] ^ d[55] ^ d[54] ^ d[53] ^ d[52] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[44] ^ d[43] ^ d[42] ^ d[41] ^ d[39] ^ d[38] ^ d[36] ^ d[32] ^ d[31] ^ d[30] ^ d[26] ^ d[25] ^ d[24] ^ d[23] ^ d[22] ^ d[21] ^ d[20] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[12] ^ d[10] ^ d[7] ^ d[6] ^ d[5] ^ d[2] ^ d[1] ^ c[1] ^ c[2] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[14] ^ c[15] ^ c[17] ^ c[18] ^ c[20] ^ c[21];
    crcf0 = newcrc;
  end
  endfunction

//synthesis translate_off
function [7:0] degree;
   input [255:0]  data;
   reg   [7:0]    i;
   begin
      i=8'b0;
      while((data>>1)>0)
      begin
         data=(data>>1);
         i=i+8'b1;
      end
      degree=i;
   end
endfunction

function    [23:0]      crc_func_0;
   input    [255:0]     data;
   reg      [255:0]     poly;
   reg      [7:0]       dataDegree;
   reg      [7:0]       polDegree;
   begin
      poly = {{233'h0},{23'h5d6dcb}};
      polDegree=degree(poly);
      data=(data<<polDegree);
      dataDegree=degree(data);
      while(dataDegree > polDegree)
      begin
         poly = {{233'h0},{23'h5D6DCB}};
         poly=(poly<<(dataDegree-polDegree));
         data=(data^poly);
         dataDegree=degree(data);
      end
      crc_func_0=data[23:0];
   end
endfunction

function    [23:0]      crc_func_1;
   input    [255:0]     data;
   reg      [255:0]     poly;
   reg      [7:0]       dataDegree;
   reg      [7:0]       polDegree;
   begin
      poly = {{232'h0},{24'h864cfb}};
      polDegree=degree(poly);
      data=(data<<polDegree);
      dataDegree=degree(data);
      while(dataDegree > polDegree)
      begin
         poly = {{232'h0},{24'h864cfb}};
         poly=(poly<<(dataDegree-polDegree));
         data=(data^poly);
         dataDegree=degree(data);
      end
      crc_func_1=data[23:0];
   end
endfunction

function [63:0] timestamp;
   input [31:0]  counter;   
   input [31:0]  carry_out;
   begin
      timestamp = ((carry_out)*(2**32-1) + counter)*TIMECLK;

   end
endfunction
//synthesis translate_on

   //--------------------- Internal Parameter-------------------------
   localparam NUM_STATES = 15;

   localparam SKIP_HDR    = 1;
   localparam WORD2_CHECK_IPV4    = 2;
   localparam WORD3_CHECK_TCP    = 4;
   localparam WORD4_IP_ADDR    = 8;
   localparam WORD5_TCP_PORT    = 16;
   localparam WORD6_TCP_ACK    = 32;
   localparam HASH_FOR_ACK    = 64;
   localparam HASH_FOR_DATA    = 128;
   localparam TEMP    = 256;
   localparam RECORD    = 512;
   localparam QUERYTEMP    = 1024;
   localparam QUERY    = 2048;
   localparam TUPLE_FOR_ACK    = 4096;
   localparam TUPLE_FOR_DATA    = 8192;
   localparam PAYLOAD            = 16384;
   
   localparam TIMECLK         = 1/(125*10**6);
   localparam TIMER_LIMIT      = 32'hffff_ffff;

   localparam ICMP        = 'h01;
   localparam TCP        = 'h06;
   localparam UDP        = 'h11;
   localparam SCTP        = 'h84;
   //------------------------- Signals-------------------------------

   wire [DATA_WIDTH-1:0]         in_fifo_data_dout;
   wire [CTRL_WIDTH-1:0]         in_fifo_ctrl_dout;

   wire [DATA_WIDTH-1:0]         pacote_data_dout;
   wire [CTRL_WIDTH-1:0]         pacote_ctrl_dout;

   wire                          in_fifo_nearly_full;
   wire                          in_fifo_empty;

   wire                          pacote_nearly_full;
   wire                          pacote_empty;

   reg                           in_fifo_rd_en;
   reg                           out_wr_int;

   /*reg                           pacote_rd_en;
   reg                           pacote_wr_en;*/

   reg [NUM_STATES-1:0]          state;
   reg [NUM_STATES-1:0]          state_next;

   reg[255:0]			            tuple_next;
   reg[255:0]			            tuple;

   reg[31:0]			            seqnum_next;
   reg[31:0]			            seqnum;

   reg[31:0]			            acknum_next;
   reg[31:0]			            acknum;

   reg[31:0]			            srcip_next;
   reg[31:0]			            srcip;

   reg[31:0]			            dstip_next;
   reg[31:0]			            dstip;

   reg[15:0]			            srcport_next;
   reg[15:0]			            srcport;

   reg[15:0]			            dstport_next;
   reg[15:0]			            dstport;

   reg[15:0]			            length_next;
   reg[15:0]			            length;

   /*reg[CRC_ADDR_WIDTH-1:0]		   hash_0_next;
   reg[CRC_ADDR_WIDTH-1:0]		   hash_0;

   reg[CRC_ADDR_WIDTH-1:0]		   hash_1_next;
   reg[CRC_ADDR_WIDTH-1:0]		   hash_1;*/
   
   /*wire                          sram0_tri_en;
   wire                          sram1_tri_en;

   wire                          sram0_we;
   wire                          sram1_we;*/

   //reg[SRAM_ADDR_WIDTH-1:0]		hash_0_next;
   reg[23:0]		               hash_0_next;

   //reg[SRAM_ADDR_WIDTH-1:0]		hash_1_next;
   reg[23:0]		               hash_1_next;

   reg                           datapkt;
   reg                           datapkt_next;

   reg                           isack;
   reg                           isack_next;

   reg                            data_pkt_next;
   reg                            ack_pkt_next;

   wire [31:0]                    num_pkts_gen;
   reg [31:0]                     num_pkts;
   reg [31:0]                     num_pkts_next;

   reg [31:0]                     num_TCP_pkts;
   reg [31:0]                     num_TCP_pkts_next;
   wire [31:0]                    num_TCP_pkts_gen;

   reg [31:0]                     num_ICMP_pkts;
   reg [31:0]                     num_ICMP_pkts_next;
   wire [31:0]                    num_ICMP_pkts_gen;

   reg [31:0]                     num_SCTP_pkts;
   reg [31:0]                     num_SCTP_pkts_next;
   wire [31:0]                    num_SCTP_pkts_gen;

   reg [31:0]                     num_UDP_pkts;
   reg [31:0]                     num_UDP_pkts_next;
   wire [31:0]                    num_UDP_pkts_gen;

   reg [31:0]                     num_ACK_pkts;
   reg [31:0]                     num_ACK_pkts_next;
   wire [31:0]                    num_ACK_pkts_gen;

   reg [31:0]                     num_escrita;
   reg [31:0]                     num_escrita_next;
   wire [31:0]                    num_escrita_gen;

   reg [31:0]                     num_leitura;
   reg [31:0]                     num_leitura_next;
   wire [31:0]                    num_leitura_gen;

   wire [31:0]                    tuple_PSRC_gen;
   wire [31:0]                    tuple_PDST_gen;
   wire [31:0]                    tuple_IPSRC_gen;
   wire [31:0]                    tuple_IPDST_gen;
   wire [31:0]                    tuple_ACKNUM_gen;
   
   //reg                            wr_0_req_aux;

   /*reg                           ctrl_flag;
   reg                           ctrl_flag_next;*/
   //------------------------- Local assignments -------------------------------

   assign in_rdy     = !in_fifo_nearly_full;
   assign out_wr     = out_wr_int;
   assign num_pkts_gen = num_pkts;
   assign num_TCP_pkts_gen = num_TCP_pkts;
   assign num_SCTP_pkts_gen = num_SCTP_pkts;
   assign num_UDP_pkts_gen = num_UDP_pkts;
   assign num_ICMP_pkts_gen = num_ICMP_pkts;
   assign num_ACK_pkts_gen = num_ACK_pkts;
   assign num_escrita_gen = num_escrita;
   assign num_leitura_gen = num_leitura;

   assign tuple_PSRC_gen = tuple[15:0];
   assign tuple_PDST_gen = tuple[31:16];
   assign tuple_IPSRC_gen = tuple[63:32];
   assign tuple_IPDST_gen = tuple[95:64];
   assign tuple_ACKNUM_gen = tuple[127:96];

   fallthrough_small_fifo #(
      .WIDTH(CTRL_WIDTH+DATA_WIDTH),
      .MAX_DEPTH_BITS(3)
   ) input_fifo (
      .din           ({in_ctrl, in_data}),   // Data in
      .wr_en         (in_wr),                // Write enable
      .rd_en         (in_fifo_rd_en),        // Read the next word
      .dout          ({in_fifo_ctrl_dout, in_fifo_data_dout}),
      .full          (),
      .nearly_full   (in_fifo_nearly_full),
      .prog_full     (),
      .empty         (in_fifo_empty),
      .reset         (reset),
      .clk           (clk)
   );

   generic_regs
   #(
      .UDP_REG_SRC_WIDTH   (UDP_REG_SRC_WIDTH),
      .TAG                 (`SIMULACAO_BLOCK_ADDR),                 // Tag -- eg. MODULE_TAG
      .REG_ADDR_WIDTH      (`SIMULACAO_REG_ADDR_WIDTH),                 // Width of block addresses -- eg. MODULE_REG_ADDR_WIDTH
      .NUM_COUNTERS        (0),                 // Number of counters
      .NUM_SOFTWARE_REGS   (0),                 // Number of sw regs
      .NUM_HARDWARE_REGS   (12)                  // Number of hw regs
   ) module_regs (
      .reg_req_in       (reg_req_in),
      .reg_ack_in       (reg_ack_in),
      .reg_rd_wr_L_in   (reg_rd_wr_L_in),
      .reg_addr_in      (reg_addr_in),
      .reg_data_in      (reg_data_in),
      .reg_src_in       (reg_src_in),

      .reg_req_out      (reg_req_out),
      .reg_ack_out      (reg_ack_out),
      .reg_rd_wr_L_out  (reg_rd_wr_L_out),
      .reg_addr_out     (reg_addr_out),
      .reg_data_out     (reg_data_out),
      .reg_src_out      (reg_src_out),

      // --- counters interface
      .counter_updates  (),
      .counter_decrement(),

      // --- SW regs interface
      .software_regs    (),

      // --- HW regs interface
      .hardware_regs    ({num_pkts_gen,num_TCP_pkts_gen,num_UDP_pkts_gen,num_ICMP_pkts_gen,num_ACK_pkts_gen,num_escrita_gen,num_leitura_gen,tuple_ACKNUM_gen,tuple_IPDST_gen,tuple_IPSRC_gen,tuple_PDST_gen,tuple_PSRC_gen}),

      .clk              (clk),
      .reset            (reset)
    );

   //------------------------- Logic-------------------------------

   always @(*) begin
      out_ctrl = in_fifo_ctrl_dout;
      out_data = in_fifo_data_dout;
      ////////////////////////////
      state_next = state;
      tuple_next = tuple;
      hash_0_next = hash_0;
      hash_1_next = hash_1;

      seqnum_next = seqnum;
      acknum_next = acknum;
      srcip_next = srcip;
      dstip_next = dstip;
      srcport_next = srcport;
      dstport_next = dstport;

      datapkt_next = datapkt;
      isack_next = isack;
      length_next = length;
      //////////////////////////// colocar if ("in_fifo_empty ...
      in_fifo_rd_en = 0; // = (!in_fifo_empty && out_rdy)
      out_wr_int = 0;

      data_pkt_next = data_pkt;
      ack_pkt_next = ack_pkt;
      num_pkts_next = num_pkts;
      num_ACK_pkts_next = num_ACK_pkts;
      num_TCP_pkts_next = num_TCP_pkts;
      num_ICMP_pkts_next = num_ICMP_pkts;
      num_UDP_pkts_next = num_UDP_pkts;
      num_SCTP_pkts_next = num_SCTP_pkts;
      num_escrita_next = num_escrita;
      num_leitura_next = num_leitura;
      
      case(state)
         // Espera por CTRL == 0 (Inicio do pacote)
         SKIP_HDR: begin
         // Wait for data to be in the FIFO and the output to be ready
         // Espera por dado na FIFO e proximo modulo estiver pronto para ler 
            //$display("SKIP HDR\n");
            if (!in_fifo_empty && out_rdy) begin
               out_wr_int = 1;
               in_fifo_rd_en = 1;
			      if(in_fifo_ctrl_dout == 'h0) begin
				      state_next = WORD2_CHECK_IPV4;
                  num_pkts_next = num_pkts_next+1;
                  //$display("numero de pacotes: %h\n",num_pkts_next);
                  //ctrl_flag_next = 1;
			      end
		      end
	      end //SKIP_HEADER
         WORD2_CHECK_IPV4: begin
            //$display("WORD2\n");
		      if (!in_fifo_empty && out_rdy) begin
           	   out_wr_int = 1;
           	   in_fifo_rd_en = 1;
			      if(in_fifo_data_dout[15:12] != 4'h4) 
                  state_next = PAYLOAD;
               else begin
                  //$display("ack0 %h ack1 %h\n",wr_0_ack, wr_1_ack);
                  state_next = WORD3_CHECK_TCP;
               end
            end
         end 
         WORD3_CHECK_TCP: begin
            //$display("WORD3\n");
            if (!in_fifo_empty && out_rdy) begin
           	   out_wr_int = 1;
           	   in_fifo_rd_en = 1;
               case(in_fifo_data_dout[7:0]) //protocolo
                  ICMP: begin
                     num_ICMP_pkts_next = num_ICMP_pkts_next + 1;
                     //$display("TCP:%03d, UDP: %03d, ICMP: %03d, SCTP %03d\n", num_TCP_pkts_next,num_UDP_pkts_next,num_ICMP_pkts_next,num_SCTP_pkts_next);
                     state_next = PAYLOAD;
                  end
                  TCP: begin
                     num_TCP_pkts_next = num_TCP_pkts_next + 1;
                     $display("TCP: %03d, UDP: %03d, ICMP: %03d, SCTP: %03d\n", num_TCP_pkts_next,num_UDP_pkts_next,num_ICMP_pkts_next,num_SCTP_pkts_next);
                     //$display("TCP: %x, UDP: %x, ICMP: %x, SCTP: %x\n", num_TCP_pkts_next,num_UDP_pkts_next,num_ICMP_pkts_next,num_SCTP_pkts_next);
                     length_next=in_fifo_data_dout[63:48]; //total_length
                     state_next = WORD4_IP_ADDR;
                  end
                  UDP: begin
                     num_UDP_pkts_next = num_UDP_pkts_next + 1;
                     //$display("TCP: %03d, UDP: %03d, ICMP: %03d, SCTP: %03d\n", num_TCP_pkts_next,num_UDP_pkts_next,num_ICMP_pkts_next,num_SCTP_pkts_next);
                     //$display("TCP: %x, UDP: %x, ICMP: %x, SCTP: %x\n", num_TCP_pkts_next,num_UDP_pkts_next,num_ICMP_pkts_next,num_SCTP_pkts_next);
                     state_next = PAYLOAD;
                  end
                  SCTP: begin
                     num_SCTP_pkts_next = num_SCTP_pkts_next + 1;
                     //$display("TCP:%03d, UDP: %03d, ICMP: %03d, SCTP: %03d\n", num_TCP_pkts_next,num_UDP_pkts_next,num_ICMP_pkts_next,num_SCTP_pkts_next);
                     //$display("TCP: %x, UDP: %x, ICMP: %x, SCTP: %x\n", num_TCP_pkts_next,num_UDP_pkts_next,num_ICMP_pkts_next,num_SCTP_pkts_next);
                     state_next = PAYLOAD;
                  end
                  default: begin
                     state_next = PAYLOAD;
                  end
               endcase
			      /*if(in_fifo_data_dout[7:0] != 8'h6) begin
                  state_next = PAYLOAD;
               end else begin
                  length_next=in_fifo_data_dout[63:48]; //total_length
                  state_next = WORD4_IP_ADDR;
               end*/
            end
         end 
         WORD4_IP_ADDR: begin
            //$display("WORD4\n");
            if (!in_fifo_empty && out_rdy) begin
           	   out_wr_int = 1;
           	   in_fifo_rd_en = 1;
               srcip_next = in_fifo_data_dout[47:16]; //srcIP
//hash_0_next = crcf0({(256-129){tuple[255:129]},(1){'b0},(129-96){seqnum},(96){tuple[95:0]}}, 256'h0);
               dstip_next[31:16] = {in_fifo_data_dout[15:0]}; //dstIp1
               state_next = WORD5_TCP_PORT;
            end
         end  
         WORD5_TCP_PORT: begin
            //$display("WORD5\n");
            if (!in_fifo_empty && out_rdy) begin
           	   out_wr_int = 1;
           	   in_fifo_rd_en = 1;
               //tuple[15:0]=in_fifo_data_dout[47:32]; //SRC_PORT
               //tuple[31:16]=in_fifo_data_dout[31:16]; //DST_PORT
               //tuple_next[31:0]=in_fifo_data_dout[47:16]; //SRC+DST PORT
               //tuple_next[47:32]=in_fifo_data_dout[63:48]; //DST_IP PART II
               dstip_next[15:0] = in_fifo_data_dout[63:48]; //dstIp2
               srcport_next = in_fifo_data_dout[47:32]; //srcPort
               dstport_next = in_fifo_data_dout[31:16]; //dstPort
               seqnum_next[31:16] = in_fifo_data_dout[15:0]; //SEQ PART I
               state_next = WORD6_TCP_ACK;
            end
         end 
         WORD6_TCP_ACK: begin
            //$display("WORD6\n");
            if (!in_fifo_empty && out_rdy) begin
           	   out_wr_int = 1;
           	   in_fifo_rd_en = 1;
               seqnum_next[15:0] = in_fifo_data_dout[63:48]; //SEQ PART II
               acknum_next = in_fifo_data_dout[47:16];
               if(in_fifo_data_dout[4]) begin //ACK flag
                  //$display("packet ack send\n");
                  isack_next = 'b1;
                  num_ACK_pkts_next = num_ACK_pkts_next + 1;
                  state_next = TUPLE_FOR_ACK;
                  //tuple_next[128:96]={(128-96){in_fifo_data_dout[63:48]}}; //seq
               end
               else begin//pkt is not ack
                  datapkt_next = 1;
                  state_next = TUPLE_FOR_DATA;
               end
               //state_next = WORD7_HASH;
            end
         end
//before alteration, out_wr_int and in_fifo_rd_en was in 0 up to PAYLOAD
         TUPLE_FOR_ACK:  begin
            $display("TUPLEACK\n");
            if (!in_fifo_empty && out_rdy) begin
           	   out_wr_int = 0;
           	   in_fifo_rd_en = 0;
               //inv{IDFlow}: src<>dst
               tuple_next[15:0]={(16){dstport}};
               tuple_next[31:16]={(16){srcport}};
               tuple_next[63:32]={(32){dstip}};
               tuple_next[95:64]={(32){srcip}};
               tuple_next[127:96]={(32){acknum}};
               tuple_next[255:128]={(256-128){1'b0}};

               state_next = HASH_FOR_ACK;
            end
         end
         TUPLE_FOR_DATA:  begin
            $display("TUPLEDATA\n");
            if (!in_fifo_empty && out_rdy) begin
           	   out_wr_int = 0;
           	   in_fifo_rd_en = 0;
               //{IDFlow}: dst<>src, sequence=seq+length+1
               //tuple_next={{128'b0},(32){seqnum+length+1},(32){dstip},(32){srcip},(16){dstport},(16){srcport}};
               tuple_next[15:0]={(16){srcport}};
               tuple_next[31:16]={(16){dstport}};
               tuple_next[63:32]={(32){srcip}};
               tuple_next[95:64]={(32){dstip}};
               tuple_next[127:96]={(32){seqnum+length+1}};
               tuple_next[255:128]={(256-128){1'b0}};

               state_next = HASH_FOR_DATA;
            end
         end
         HASH_FOR_ACK:  begin
            $display("HASHACK\n");
            if (!in_fifo_empty && out_rdy) begin
               $display("ACK tuple: %h\n",tuple[127:0]);
           	   out_wr_int = 0;
           	   in_fifo_rd_en = 0;
               hash_0_next = {2'b0,crcf0(tuple, 256'h0)};
               hash_1_next = {1'b0,crcf1(tuple, 256'h0)}; 
               state_next = TEMP;
               ack_pkt_next = 1'b1;
               //ack_pkt = 1'b1;
            end
         end
         HASH_FOR_DATA:  begin
            $display("HASHDATA\n");
            if (!in_fifo_empty && out_rdy) begin
               $display("DATA tuple: %h\n",tuple[127:0]);
           	   out_wr_int = 0;
           	   in_fifo_rd_en = 0;
               hash_0_next = crcf0(tuple, 256'h0);
               hash_1_next = crcf1(tuple, 256'h0);
               state_next = TEMP;
               data_pkt_next = 1'b1;
            end
         end
         TEMP:  begin
            $display("TEMP\n");
            {data_pkt_next,ack_pkt_next} = 2'b0;
            if (!in_fifo_empty && out_rdy) begin
                  out_wr_int = 0;
                  in_fifo_rd_en = 0;
               if(data_proc||ack_proc) begin
                  $display("dataproc: %x\n", hash_0_next);
                  //{data_pkt_next,ack_pkt_next} = 2'b0;
                  //{data_pkt,ack_pkt} = 2'b0;
 //if packet is ack and data, after reading must be write operation
                  if(length > 0 && isack) begin
                     datapkt_next = 0;
                     isack_next = 0;
                     state_next = TUPLE_FOR_DATA;
                  end
                  else
                     state_next = PAYLOAD;
               end
               else 
                  state_next = TEMP;
            end
         end
		   PAYLOAD: begin
            $display("PAYLOAD\n");
		      if (!in_fifo_empty && out_rdy) begin
           	   out_wr_int = 1;
           	   in_fifo_rd_en = 1;
               hash_0_next = 0;
               hash_1_next = 0;
			      //CHECA POR FIM DO PACOTE
		   	   if(in_fifo_ctrl_dout != 'h0)
				      state_next = SKIP_HDR;
               else
				      state_next = PAYLOAD;
		      end
	      end //PAYLOAD
	   endcase //case(state)
   end //always

   always @(posedge clk) begin
	   if(reset) begin
      ////////////////////-Sram
         {data_pkt,ack_pkt} <= 2'b0;
      ////////////////////-Sram
		   state <= SKIP_HDR;
         tuple <= 256'h0;
         seqnum <= 32'h0;
         acknum <= 32'h0;
         hash_0 <= {{SRAM_ADDR_WIDTH}{1'b0}};
         hash_1 <= {{SRAM_ADDR_WIDTH}{1'b0}}; //24'h0;

         srcip <=32'h0;
         dstip <=32'h0;
         srcport <=16'h0;
         dstport <=16'h0;

         isack <= 0;
         datapkt <= 0;
         length <= 0;

         num_pkts <= 0;
         num_UDP_pkts <= 0;
         num_SCTP_pkts <= 0;
         num_ICMP_pkts <= 0;
         num_TCP_pkts <= 0;
         num_ACK_pkts <= 0;
         num_escrita <= 0;
         num_leitura <= 0;
	   end
	   else begin
         //if(state_next != SKIP_HDR) begin
            //$display("state_next: %d\n", 30'h3fff_ffff);
            //$display("fifo_data_dout: %h\n", in_fifo_data_dout);
            //$display("hash_0: %h, hash_1: %h\n", hash_0_next, hash_1_next);
         //end
         /////////////////--Sram
         //if(state_next == WORD4_IP_ADDR) begin
            //wr_0_req_aux <= 0;
            //$display("length: %d, %x\n", length_next,length_next);
         //end
         //else if(state_next == WORD5_TCP_PORT) begin
            //$display("src ip: %03d.%03d.%03d.%03d\n", srcip_next[31:24],srcip_next[23:16],srcip_next[15:8],srcip_next[7:0]);
         //end
         //else if(state_next == WORD6_TCP_ACK) begin
            //$display("dst ip: %03d.%03d.%03d.%03d\n", dstip_next[31:24],dstip_next[23:16],dstip_next[15:8],dstip_next[7:0]);
            //$display("dst port: %d, %x\n",dstport_next,dstport_next);
            //$display("src port: %d, %x\n",srcport_next,srcport_next);
         //end
         if(in_fifo_nearly_full)
            $display("in_fifo_nearly_full: %d\n",in_fifo_nearly_full);
         data_pkt <= data_pkt_next;
         ack_pkt <= ack_pkt_next;
		   state <= state_next;
         tuple <= tuple_next;

         seqnum <= seqnum_next;
         acknum <= acknum_next;
         srcip <= srcip_next;
         dstip <= dstip_next;
         srcport <= srcport_next;
         dstport <= dstport_next;

         hash_0 <= hash_0_next;
         hash_1 <= hash_1_next;
         isack <= isack_next;
         datapkt <= datapkt_next;
         length <= length_next;
         num_pkts <= num_pkts_next;
         num_TCP_pkts <= num_TCP_pkts_next;

         num_ICMP_pkts <= num_ICMP_pkts_next;
         num_UDP_pkts <= num_UDP_pkts_next;
         num_SCTP_pkts <= num_SCTP_pkts_next;
         num_ACK_pkts <= num_ACK_pkts_next;
         num_escrita <= num_escrita_next;
         num_leitura <= num_leitura_next;
	   end
   end
endmodule
